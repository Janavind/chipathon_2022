magic
tech sky130B
magscale 1 2
timestamp 1669671049
<< viali >>
rect 4721 47209 4755 47243
rect 5365 47209 5399 47243
rect 6009 47209 6043 47243
rect 7113 47209 7147 47243
rect 7757 47209 7791 47243
rect 8401 47209 8435 47243
rect 9137 47209 9171 47243
rect 10241 47209 10275 47243
rect 11161 47209 11195 47243
rect 12449 47209 12483 47243
rect 13553 47209 13587 47243
rect 15025 47209 15059 47243
rect 20637 47209 20671 47243
rect 24041 47209 24075 47243
rect 26065 47209 26099 47243
rect 43913 47209 43947 47243
rect 45201 47209 45235 47243
rect 46489 47209 46523 47243
rect 38209 47141 38243 47175
rect 38945 47141 38979 47175
rect 41429 47141 41463 47175
rect 44557 47141 44591 47175
rect 15669 47073 15703 47107
rect 19441 47073 19475 47107
rect 19993 47073 20027 47107
rect 22569 47073 22603 47107
rect 24593 47073 24627 47107
rect 29745 47073 29779 47107
rect 31217 47073 31251 47107
rect 33241 47073 33275 47107
rect 16313 47005 16347 47039
rect 17509 47005 17543 47039
rect 18429 47005 18463 47039
rect 18521 47005 18555 47039
rect 19901 47005 19935 47039
rect 20453 47005 20487 47039
rect 21465 47005 21499 47039
rect 22017 47005 22051 47039
rect 22109 47005 22143 47039
rect 23397 47005 23431 47039
rect 25145 47005 25179 47039
rect 25421 47005 25455 47039
rect 25605 47005 25639 47039
rect 27721 47005 27755 47039
rect 27997 47005 28031 47039
rect 28181 47005 28215 47039
rect 28917 47005 28951 47039
rect 30757 47005 30791 47039
rect 31125 47005 31159 47039
rect 33517 47005 33551 47039
rect 33701 47005 33735 47039
rect 34161 47005 34195 47039
rect 35357 47005 35391 47039
rect 35541 47005 35575 47039
rect 35725 47005 35759 47039
rect 36369 47005 36403 47039
rect 37473 47005 37507 47039
rect 38393 47005 38427 47039
rect 39129 47005 39163 47039
rect 40877 47005 40911 47039
rect 41613 47005 41647 47039
rect 42625 47005 42659 47039
rect 43269 47005 43303 47039
rect 45845 47005 45879 47039
rect 17969 46937 18003 46971
rect 27169 46937 27203 46971
rect 30297 46937 30331 46971
rect 32689 46937 32723 46971
rect 34897 46937 34931 46971
rect 17325 46869 17359 46903
rect 21281 46869 21315 46903
rect 29101 46869 29135 46903
rect 40601 46869 40635 46903
rect 16129 46665 16163 46699
rect 25881 46597 25915 46631
rect 27813 46597 27847 46631
rect 33701 46597 33735 46631
rect 41981 46597 42015 46631
rect 6929 46529 6963 46563
rect 14657 46529 14691 46563
rect 15577 46529 15611 46563
rect 16313 46529 16347 46563
rect 17233 46529 17267 46563
rect 17693 46529 17727 46563
rect 18245 46529 18279 46563
rect 18429 46529 18463 46563
rect 18981 46529 19015 46563
rect 19165 46529 19199 46563
rect 20177 46529 20211 46563
rect 21373 46529 21407 46563
rect 22109 46529 22143 46563
rect 22845 46529 22879 46563
rect 23480 46529 23514 46563
rect 23673 46529 23707 46563
rect 24041 46529 24075 46563
rect 24133 46529 24167 46563
rect 24317 46529 24351 46563
rect 26249 46529 26283 46563
rect 26341 46529 26375 46563
rect 29101 46529 29135 46563
rect 29653 46529 29687 46563
rect 30481 46529 30515 46563
rect 31309 46529 31343 46563
rect 33057 46529 33091 46563
rect 33241 46529 33275 46563
rect 34161 46529 34195 46563
rect 34437 46529 34471 46563
rect 34621 46529 34655 46563
rect 35173 46529 35207 46563
rect 35633 46529 35667 46563
rect 36461 46529 36495 46563
rect 38301 46529 38335 46563
rect 38485 46529 38519 46563
rect 39589 46529 39623 46563
rect 40233 46529 40267 46563
rect 43269 46529 43303 46563
rect 44557 46529 44591 46563
rect 45201 46529 45235 46563
rect 45845 46529 45879 46563
rect 17785 46461 17819 46495
rect 20913 46461 20947 46495
rect 21469 46461 21503 46495
rect 26433 46461 26467 46495
rect 27169 46461 27203 46495
rect 31125 46461 31159 46495
rect 32781 46461 32815 46495
rect 34805 46461 34839 46495
rect 36185 46461 36219 46495
rect 36645 46461 36679 46495
rect 37473 46461 37507 46495
rect 38025 46461 38059 46495
rect 39497 46461 39531 46495
rect 40693 46461 40727 46495
rect 43913 46461 43947 46495
rect 22293 46393 22327 46427
rect 25421 46393 25455 46427
rect 30297 46393 30331 46427
rect 41337 46393 41371 46427
rect 42625 46393 42659 46427
rect 19441 46325 19475 46359
rect 20361 46325 20395 46359
rect 24961 46325 24995 46359
rect 16957 46121 16991 46155
rect 18705 46121 18739 46155
rect 19533 46121 19567 46155
rect 27261 46121 27295 46155
rect 30205 46121 30239 46155
rect 36369 46121 36403 46155
rect 42349 46121 42383 46155
rect 43637 46121 43671 46155
rect 44281 46121 44315 46155
rect 31677 46053 31711 46087
rect 42993 46053 43027 46087
rect 18061 45985 18095 46019
rect 21465 45985 21499 46019
rect 22385 45985 22419 46019
rect 23397 45985 23431 46019
rect 33057 45985 33091 46019
rect 35541 45985 35575 46019
rect 36829 45985 36863 46019
rect 39221 45985 39255 46019
rect 40601 45985 40635 46019
rect 16313 45917 16347 45951
rect 17417 45917 17451 45951
rect 17509 45917 17543 45951
rect 17969 45917 18003 45951
rect 18889 45917 18923 45951
rect 19993 45917 20027 45951
rect 20105 45917 20139 45951
rect 21741 45917 21775 45951
rect 21837 45917 21871 45951
rect 22477 45917 22511 45951
rect 23305 45917 23339 45951
rect 23581 45917 23615 45951
rect 25053 45917 25087 45951
rect 25421 45917 25455 45951
rect 25513 45917 25547 45951
rect 26249 45917 26283 45951
rect 26341 45917 26375 45951
rect 26801 45917 26835 45951
rect 26985 45917 27019 45951
rect 28917 45917 28951 45951
rect 29193 45917 29227 45951
rect 29745 45917 29779 45951
rect 30113 45917 30147 45951
rect 30941 45917 30975 45951
rect 32045 45917 32079 45951
rect 32689 45917 32723 45951
rect 33885 45917 33919 45951
rect 34897 45917 34931 45951
rect 36921 45917 36955 45951
rect 37289 45917 37323 45951
rect 37473 45917 37507 45951
rect 38301 45917 38335 45951
rect 39129 45917 39163 45951
rect 40693 45917 40727 45951
rect 41153 45917 41187 45951
rect 41245 45917 41279 45951
rect 20545 45849 20579 45883
rect 24593 45849 24627 45883
rect 28457 45849 28491 45883
rect 29009 45849 29043 45883
rect 33517 45849 33551 45883
rect 34069 45849 34103 45883
rect 38393 45849 38427 45883
rect 27905 45781 27939 45815
rect 41705 45781 41739 45815
rect 23673 45577 23707 45611
rect 24869 45509 24903 45543
rect 34713 45509 34747 45543
rect 35725 45509 35759 45543
rect 40693 45509 40727 45543
rect 17877 45441 17911 45475
rect 18797 45441 18831 45475
rect 18981 45441 19015 45475
rect 19349 45441 19383 45475
rect 20545 45441 20579 45475
rect 20913 45441 20947 45475
rect 21097 45441 21131 45475
rect 22477 45441 22511 45475
rect 22845 45441 22879 45475
rect 23213 45441 23247 45475
rect 25513 45441 25547 45475
rect 25881 45441 25915 45475
rect 26065 45441 26099 45475
rect 26525 45441 26559 45475
rect 28181 45441 28215 45475
rect 28549 45441 28583 45475
rect 28641 45441 28675 45475
rect 29377 45441 29411 45475
rect 30113 45441 30147 45475
rect 31033 45441 31067 45475
rect 31493 45441 31527 45475
rect 33333 45441 33367 45475
rect 33701 45441 33735 45475
rect 35081 45441 35115 45475
rect 35265 45441 35299 45475
rect 36461 45441 36495 45475
rect 36737 45441 36771 45475
rect 38117 45441 38151 45475
rect 38485 45441 38519 45475
rect 39129 45441 39163 45475
rect 40325 45441 40359 45475
rect 40785 45441 40819 45475
rect 41521 45441 41555 45475
rect 42625 45441 42659 45475
rect 18337 45373 18371 45407
rect 19257 45373 19291 45407
rect 22937 45373 22971 45407
rect 23121 45373 23155 45407
rect 25605 45373 25639 45407
rect 29285 45373 29319 45407
rect 30205 45373 30239 45407
rect 34069 45373 34103 45407
rect 36277 45373 36311 45407
rect 36921 45373 36955 45407
rect 38577 45373 38611 45407
rect 40601 45373 40635 45407
rect 43821 45373 43855 45407
rect 17233 45305 17267 45339
rect 27997 45305 28031 45339
rect 30849 45305 30883 45339
rect 37933 45305 37967 45339
rect 39865 45305 39899 45339
rect 20085 45237 20119 45271
rect 24409 45237 24443 45271
rect 27261 45237 27295 45271
rect 39313 45237 39347 45271
rect 43269 45237 43303 45271
rect 18337 45033 18371 45067
rect 24041 45033 24075 45067
rect 34161 45033 34195 45067
rect 40049 45033 40083 45067
rect 42257 45033 42291 45067
rect 24869 44965 24903 44999
rect 28733 44965 28767 44999
rect 30021 44965 30055 44999
rect 31125 44965 31159 44999
rect 35173 44965 35207 44999
rect 20637 44897 20671 44931
rect 23397 44897 23431 44931
rect 25421 44897 25455 44931
rect 28089 44897 28123 44931
rect 37013 44897 37047 44931
rect 40693 44897 40727 44931
rect 41245 44897 41279 44931
rect 42717 44897 42751 44931
rect 18153 44829 18187 44863
rect 19993 44829 20027 44863
rect 20545 44829 20579 44863
rect 22017 44829 22051 44863
rect 22937 44829 22971 44863
rect 23213 44829 23247 44863
rect 24685 44829 24719 44863
rect 25973 44829 26007 44863
rect 26249 44829 26283 44863
rect 26433 44829 26467 44863
rect 27629 44829 27663 44863
rect 27997 44829 28031 44863
rect 28917 44829 28951 44863
rect 29745 44829 29779 44863
rect 30389 44829 30423 44863
rect 31953 44829 31987 44863
rect 32045 44829 32079 44863
rect 32321 44829 32355 44863
rect 33609 44829 33643 44863
rect 33701 44829 33735 44863
rect 34897 44829 34931 44863
rect 35541 44829 35575 44863
rect 35725 44829 35759 44863
rect 37289 44829 37323 44863
rect 37473 44829 37507 44863
rect 38209 44829 38243 44863
rect 38669 44829 38703 44863
rect 38945 44829 38979 44863
rect 39313 44829 39347 44863
rect 41521 44829 41555 44863
rect 41705 44829 41739 44863
rect 22201 44761 22235 44795
rect 27169 44761 27203 44795
rect 31585 44761 31619 44795
rect 33149 44761 33183 44795
rect 36461 44761 36495 44795
rect 19809 44693 19843 44727
rect 21925 44693 21959 44727
rect 43269 44693 43303 44727
rect 19625 44489 19659 44523
rect 21281 44489 21315 44523
rect 26341 44489 26375 44523
rect 41889 44489 41923 44523
rect 42625 44489 42659 44523
rect 18337 44421 18371 44455
rect 22845 44421 22879 44455
rect 23765 44421 23799 44455
rect 28181 44421 28215 44455
rect 33425 44421 33459 44455
rect 34989 44421 35023 44455
rect 41429 44421 41463 44455
rect 19073 44353 19107 44387
rect 19809 44353 19843 44387
rect 20361 44353 20395 44387
rect 20545 44353 20579 44387
rect 21097 44353 21131 44387
rect 22477 44353 22511 44387
rect 22937 44353 22971 44387
rect 24317 44353 24351 44387
rect 24593 44353 24627 44387
rect 24777 44353 24811 44387
rect 25237 44353 25271 44387
rect 25421 44353 25455 44387
rect 26341 44353 26375 44387
rect 27445 44353 27479 44387
rect 27813 44353 27847 44387
rect 28733 44353 28767 44387
rect 29469 44353 29503 44387
rect 29837 44353 29871 44387
rect 31217 44353 31251 44387
rect 31585 44353 31619 44387
rect 32413 44353 32447 44387
rect 34345 44353 34379 44387
rect 34529 44353 34563 44387
rect 35633 44353 35667 44387
rect 36185 44353 36219 44387
rect 37473 44353 37507 44387
rect 37933 44353 37967 44387
rect 38117 44353 38151 44387
rect 38301 44353 38335 44387
rect 38945 44353 38979 44387
rect 39313 44353 39347 44387
rect 40509 44353 40543 44387
rect 40877 44353 40911 44387
rect 22017 44285 22051 44319
rect 23121 44285 23155 44319
rect 25789 44285 25823 44319
rect 29009 44285 29043 44319
rect 30941 44285 30975 44319
rect 32781 44285 32815 44319
rect 32873 44285 32907 44319
rect 36369 44285 36403 44319
rect 40141 44285 40175 44319
rect 31493 44217 31527 44251
rect 35633 44217 35667 44251
rect 34253 44149 34287 44183
rect 39405 44149 39439 44183
rect 24041 43945 24075 43979
rect 28917 43945 28951 43979
rect 30113 43945 30147 43979
rect 31125 43945 31159 43979
rect 33241 43945 33275 43979
rect 37289 43945 37323 43979
rect 38393 43945 38427 43979
rect 40601 43945 40635 43979
rect 41797 43945 41831 43979
rect 22017 43877 22051 43911
rect 20177 43809 20211 43843
rect 26985 43809 27019 43843
rect 33701 43809 33735 43843
rect 38853 43809 38887 43843
rect 39313 43809 39347 43843
rect 40049 43809 40083 43843
rect 20545 43741 20579 43775
rect 20729 43741 20763 43775
rect 21465 43741 21499 43775
rect 21741 43741 21775 43775
rect 22293 43741 22327 43775
rect 22845 43741 22879 43775
rect 25513 43741 25547 43775
rect 26433 43741 26467 43775
rect 27445 43741 27479 43775
rect 27629 43741 27663 43775
rect 27813 43741 27847 43775
rect 28089 43741 28123 43775
rect 28365 43741 28399 43775
rect 31585 43741 31619 43775
rect 32229 43741 32263 43775
rect 33793 43741 33827 43775
rect 34161 43741 34195 43775
rect 34345 43741 34379 43775
rect 35449 43741 35483 43775
rect 35909 43741 35943 43775
rect 38577 43741 38611 43775
rect 38669 43741 38703 43775
rect 23305 43673 23339 43707
rect 24593 43673 24627 43707
rect 19717 43605 19751 43639
rect 23029 43605 23063 43639
rect 41153 43605 41187 43639
rect 28181 43401 28215 43435
rect 37565 43401 37599 43435
rect 23029 43333 23063 43367
rect 26617 43333 26651 43367
rect 32781 43333 32815 43367
rect 38301 43333 38335 43367
rect 21281 43265 21315 43299
rect 22109 43265 22143 43299
rect 23673 43265 23707 43299
rect 24041 43265 24075 43299
rect 24225 43265 24259 43299
rect 25697 43265 25731 43299
rect 25789 43265 25823 43299
rect 26157 43265 26191 43299
rect 27261 43265 27295 43299
rect 27721 43265 27755 43299
rect 28089 43265 28123 43299
rect 29929 43265 29963 43299
rect 30021 43265 30055 43299
rect 30205 43265 30239 43299
rect 33241 43265 33275 43299
rect 33609 43265 33643 43299
rect 34253 43265 34287 43299
rect 36369 43265 36403 43299
rect 36645 43265 36679 43299
rect 39405 43265 39439 43299
rect 39957 43265 39991 43299
rect 20637 43197 20671 43231
rect 22017 43197 22051 43231
rect 22569 43197 22603 43231
rect 23581 43197 23615 43231
rect 29193 43197 29227 43231
rect 29745 43197 29779 43231
rect 31401 43197 31435 43231
rect 33701 43197 33735 43231
rect 24685 43129 24719 43163
rect 30849 43129 30883 43163
rect 34989 43061 35023 43095
rect 23213 42857 23247 42891
rect 25973 42857 26007 42891
rect 31217 42789 31251 42823
rect 27445 42721 27479 42755
rect 29009 42721 29043 42755
rect 30297 42721 30331 42755
rect 30757 42721 30791 42755
rect 33149 42721 33183 42755
rect 33793 42721 33827 42755
rect 34897 42721 34931 42755
rect 35541 42721 35575 42755
rect 36461 42721 36495 42755
rect 38025 42721 38059 42755
rect 38577 42721 38611 42755
rect 39221 42721 39255 42755
rect 22661 42653 22695 42687
rect 23029 42653 23063 42687
rect 25421 42653 25455 42687
rect 25513 42653 25547 42687
rect 27077 42653 27111 42687
rect 27997 42653 28031 42687
rect 28549 42653 28583 42687
rect 30573 42653 30607 42687
rect 32413 42653 32447 42687
rect 34253 42653 34287 42687
rect 34345 42653 34379 42687
rect 37473 42653 37507 42687
rect 24961 42585 24995 42619
rect 26893 42585 26927 42619
rect 29745 42585 29779 42619
rect 28089 42517 28123 42551
rect 31769 42517 31803 42551
rect 36921 42517 36955 42551
rect 23673 42313 23707 42347
rect 26249 42313 26283 42347
rect 30113 42313 30147 42347
rect 30665 42313 30699 42347
rect 31769 42313 31803 42347
rect 32321 42313 32355 42347
rect 33885 42313 33919 42347
rect 34437 42313 34471 42347
rect 34989 42313 35023 42347
rect 36185 42313 36219 42347
rect 38117 42313 38151 42347
rect 31125 42245 31159 42279
rect 33333 42245 33367 42279
rect 36737 42245 36771 42279
rect 37473 42245 37507 42279
rect 23765 42177 23799 42211
rect 24317 42177 24351 42211
rect 25145 42177 25179 42211
rect 25513 42177 25547 42211
rect 25697 42177 25731 42211
rect 29101 42177 29135 42211
rect 29469 42177 29503 42211
rect 24593 42109 24627 42143
rect 22661 41973 22695 42007
rect 27629 41973 27663 42007
rect 35541 41973 35575 42007
rect 25053 41769 25087 41803
rect 31309 41769 31343 41803
rect 34161 41769 34195 41803
rect 34897 41701 34931 41735
rect 28917 41633 28951 41667
rect 29837 41633 29871 41667
rect 26157 41565 26191 41599
rect 26617 41565 26651 41599
rect 29929 41497 29963 41531
rect 30849 41497 30883 41531
rect 28089 41429 28123 41463
rect 24869 41225 24903 41259
rect 26525 41225 26559 41259
rect 27261 41225 27295 41259
rect 28549 41225 28583 41259
rect 29193 41225 29227 41259
rect 25513 41157 25547 41191
rect 27721 41157 27755 41191
rect 26065 41089 26099 41123
rect 29653 40885 29687 40919
rect 28825 40681 28859 40715
rect 22937 7837 22971 7871
rect 24041 7837 24075 7871
rect 24777 7837 24811 7871
rect 25605 7837 25639 7871
rect 26065 7837 26099 7871
rect 25421 7701 25455 7735
rect 21281 7497 21315 7531
rect 24869 7429 24903 7463
rect 24961 7429 24995 7463
rect 25697 7429 25731 7463
rect 22661 7361 22695 7395
rect 24685 7293 24719 7327
rect 25605 7293 25639 7327
rect 26617 7293 26651 7327
rect 22201 7157 22235 7191
rect 22937 7157 22971 7191
rect 27169 7157 27203 7191
rect 27813 7157 27847 7191
rect 24869 6953 24903 6987
rect 25697 6953 25731 6987
rect 23029 6817 23063 6851
rect 23857 6817 23891 6851
rect 27721 6817 27755 6851
rect 27997 6817 28031 6851
rect 20729 6749 20763 6783
rect 21465 6749 21499 6783
rect 22477 6749 22511 6783
rect 24593 6749 24627 6783
rect 25697 6749 25731 6783
rect 26433 6749 26467 6783
rect 23121 6681 23155 6715
rect 27813 6681 27847 6715
rect 20177 6613 20211 6647
rect 20913 6613 20947 6647
rect 21649 6613 21683 6647
rect 22293 6613 22327 6647
rect 26617 6613 26651 6647
rect 27629 6409 27663 6443
rect 20545 6341 20579 6375
rect 22569 6341 22603 6375
rect 24041 6341 24075 6375
rect 24133 6341 24167 6375
rect 25697 6341 25731 6375
rect 27629 6273 27663 6307
rect 28273 6273 28307 6307
rect 19901 6205 19935 6239
rect 20453 6205 20487 6239
rect 21097 6205 21131 6239
rect 22477 6205 22511 6239
rect 23489 6205 23523 6239
rect 24961 6205 24995 6239
rect 25605 6205 25639 6239
rect 26433 6205 26467 6239
rect 28273 6069 28307 6103
rect 29193 6069 29227 6103
rect 20821 5865 20855 5899
rect 22569 5865 22603 5899
rect 24685 5865 24719 5899
rect 25697 5865 25731 5899
rect 26433 5865 26467 5899
rect 27721 5729 27755 5763
rect 20177 5661 20211 5695
rect 20913 5661 20947 5695
rect 21649 5661 21683 5695
rect 22569 5661 22603 5695
rect 23673 5661 23707 5695
rect 24685 5661 24719 5695
rect 25421 5661 25455 5695
rect 26249 5661 26283 5695
rect 29009 5661 29043 5695
rect 22017 5593 22051 5627
rect 24041 5593 24075 5627
rect 28181 5593 28215 5627
rect 28273 5593 28307 5627
rect 29193 5593 29227 5627
rect 20085 5525 20119 5559
rect 19901 5253 19935 5287
rect 22661 5253 22695 5287
rect 24317 5253 24351 5287
rect 26617 5253 26651 5287
rect 27353 5253 27387 5287
rect 29653 5253 29687 5287
rect 29745 5253 29779 5287
rect 26525 5185 26559 5219
rect 19809 5117 19843 5151
rect 20821 5117 20855 5151
rect 22569 5117 22603 5151
rect 23213 5117 23247 5151
rect 24225 5117 24259 5151
rect 24869 5117 24903 5151
rect 27261 5117 27295 5151
rect 27629 5117 27663 5151
rect 28825 5117 28859 5151
rect 21465 5049 21499 5083
rect 19257 4981 19291 5015
rect 18245 4777 18279 4811
rect 18889 4777 18923 4811
rect 24777 4777 24811 4811
rect 27445 4777 27479 4811
rect 21189 4641 21223 4675
rect 21833 4641 21867 4675
rect 25973 4641 26007 4675
rect 28825 4641 28859 4675
rect 29101 4641 29135 4675
rect 30573 4641 30607 4675
rect 19533 4573 19567 4607
rect 20361 4573 20395 4607
rect 22845 4573 22879 4607
rect 23949 4573 23983 4607
rect 29837 4573 29871 4607
rect 21281 4505 21315 4539
rect 23213 4505 23247 4539
rect 24041 4505 24075 4539
rect 25329 4505 25363 4539
rect 25421 4505 25455 4539
rect 29009 4505 29043 4539
rect 19717 4437 19751 4471
rect 20545 4437 20579 4471
rect 29837 4437 29871 4471
rect 25421 4233 25455 4267
rect 22201 4165 22235 4199
rect 23765 4165 23799 4199
rect 28089 4165 28123 4199
rect 20361 4097 20395 4131
rect 21281 4097 21315 4131
rect 25513 4097 25547 4131
rect 26525 4097 26559 4131
rect 26617 4097 26651 4131
rect 29101 4097 29135 4131
rect 19165 4029 19199 4063
rect 22109 4029 22143 4063
rect 22385 4029 22419 4063
rect 23673 4029 23707 4063
rect 24133 4029 24167 4063
rect 27169 4029 27203 4063
rect 28181 4029 28215 4063
rect 29561 4029 29595 4063
rect 17877 3961 17911 3995
rect 19809 3961 19843 3995
rect 16129 3893 16163 3927
rect 17233 3893 17267 3927
rect 18521 3893 18555 3927
rect 20545 3893 20579 3927
rect 21373 3893 21407 3927
rect 28825 3893 28859 3927
rect 30205 3893 30239 3927
rect 18245 3689 18279 3723
rect 16313 3621 16347 3655
rect 17601 3621 17635 3655
rect 19441 3621 19475 3655
rect 31677 3621 31711 3655
rect 16957 3553 16991 3587
rect 18889 3553 18923 3587
rect 22477 3553 22511 3587
rect 22753 3553 22787 3587
rect 28549 3553 28583 3587
rect 28825 3553 28859 3587
rect 4261 3485 4295 3519
rect 5181 3485 5215 3519
rect 6009 3485 6043 3519
rect 6837 3485 6871 3519
rect 7665 3485 7699 3519
rect 8493 3485 8527 3519
rect 9321 3485 9355 3519
rect 10149 3485 10183 3519
rect 10977 3485 11011 3519
rect 11713 3485 11747 3519
rect 12357 3485 12391 3519
rect 13001 3485 13035 3519
rect 13645 3485 13679 3519
rect 15025 3485 15059 3519
rect 15669 3485 15703 3519
rect 21557 3485 21591 3519
rect 25421 3485 25455 3519
rect 26525 3485 26559 3519
rect 29745 3485 29779 3519
rect 30389 3485 30423 3519
rect 31033 3485 31067 3519
rect 32321 3485 32355 3519
rect 32965 3485 32999 3519
rect 33609 3485 33643 3519
rect 35173 3485 35207 3519
rect 35633 3485 35667 3519
rect 36277 3485 36311 3519
rect 37105 3485 37139 3519
rect 37933 3485 37967 3519
rect 39037 3485 39071 3519
rect 40417 3485 40451 3519
rect 40877 3485 40911 3519
rect 41521 3485 41555 3519
rect 42901 3485 42935 3519
rect 43361 3485 43395 3519
rect 45201 3485 45235 3519
rect 45845 3485 45879 3519
rect 46489 3485 46523 3519
rect 47133 3485 47167 3519
rect 47777 3485 47811 3519
rect 20085 3417 20119 3451
rect 20177 3417 20211 3451
rect 21097 3417 21131 3451
rect 22569 3417 22603 3451
rect 28733 3417 28767 3451
rect 21833 3349 21867 3383
rect 25421 3349 25455 3383
rect 26709 3349 26743 3383
rect 20085 3145 20119 3179
rect 22201 3077 22235 3111
rect 23857 3077 23891 3111
rect 25421 3077 25455 3111
rect 28089 3077 28123 3111
rect 29653 3077 29687 3111
rect 30297 3077 30331 3111
rect 18245 3009 18279 3043
rect 18889 3009 18923 3043
rect 20361 3009 20395 3043
rect 21373 3009 21407 3043
rect 30389 3009 30423 3043
rect 4721 2941 4755 2975
rect 7297 2941 7331 2975
rect 9229 2941 9263 2975
rect 14381 2941 14415 2975
rect 15669 2941 15703 2975
rect 17601 2941 17635 2975
rect 22109 2941 22143 2975
rect 22477 2941 22511 2975
rect 23765 2941 23799 2975
rect 24409 2941 24443 2975
rect 25329 2941 25363 2975
rect 25789 2941 25823 2975
rect 27169 2941 27203 2975
rect 28181 2941 28215 2975
rect 29377 2941 29411 2975
rect 29745 2941 29779 2975
rect 33609 2941 33643 2975
rect 39405 2941 39439 2975
rect 41337 2941 41371 2975
rect 43269 2941 43303 2975
rect 45201 2941 45235 2975
rect 4077 2873 4111 2907
rect 5365 2873 5399 2907
rect 10517 2873 10551 2907
rect 12449 2873 12483 2907
rect 13737 2873 13771 2907
rect 16313 2873 16347 2907
rect 19533 2873 19567 2907
rect 35541 2873 35575 2907
rect 2789 2805 2823 2839
rect 3433 2805 3467 2839
rect 6009 2805 6043 2839
rect 7941 2805 7975 2839
rect 8585 2805 8619 2839
rect 9873 2805 9907 2839
rect 11161 2805 11195 2839
rect 13093 2805 13127 2839
rect 15025 2805 15059 2839
rect 21373 2805 21407 2839
rect 31125 2805 31159 2839
rect 32321 2805 32355 2839
rect 32965 2805 32999 2839
rect 34253 2805 34287 2839
rect 34897 2805 34931 2839
rect 36185 2805 36219 2839
rect 37473 2805 37507 2839
rect 38117 2805 38151 2839
rect 38761 2805 38795 2839
rect 40049 2805 40083 2839
rect 40693 2805 40727 2839
rect 42625 2805 42659 2839
rect 43913 2805 43947 2839
rect 44557 2805 44591 2839
rect 45845 2805 45879 2839
rect 46489 2805 46523 2839
rect 47777 2805 47811 2839
rect 18889 2601 18923 2635
rect 21373 2601 21407 2635
rect 26433 2601 26467 2635
rect 30573 2601 30607 2635
rect 31217 2601 31251 2635
rect 5365 2533 5399 2567
rect 7941 2533 7975 2567
rect 9873 2533 9907 2567
rect 12449 2533 12483 2567
rect 17601 2533 17635 2567
rect 20637 2533 20671 2567
rect 33609 2533 33643 2567
rect 36185 2533 36219 2567
rect 40049 2533 40083 2567
rect 43913 2533 43947 2567
rect 46489 2533 46523 2567
rect 2789 2465 2823 2499
rect 7297 2465 7331 2499
rect 8585 2465 8619 2499
rect 11161 2465 11195 2499
rect 13093 2465 13127 2499
rect 15025 2465 15059 2499
rect 19993 2465 20027 2499
rect 22753 2465 22787 2499
rect 23029 2465 23063 2499
rect 24961 2465 24995 2499
rect 25513 2465 25547 2499
rect 28273 2465 28307 2499
rect 28641 2465 28675 2499
rect 32965 2465 32999 2499
rect 34897 2465 34931 2499
rect 38117 2465 38151 2499
rect 40693 2465 40727 2499
rect 42625 2465 42659 2499
rect 45201 2465 45235 2499
rect 2145 2397 2179 2431
rect 3433 2397 3467 2431
rect 4721 2397 4755 2431
rect 6009 2397 6043 2431
rect 10517 2397 10551 2431
rect 13737 2397 13771 2431
rect 15669 2397 15703 2431
rect 16313 2397 16347 2431
rect 18245 2397 18279 2431
rect 21097 2397 21131 2431
rect 22201 2397 22235 2431
rect 30113 2397 30147 2431
rect 32321 2397 32355 2431
rect 35541 2397 35575 2431
rect 37473 2397 37507 2431
rect 38761 2397 38795 2431
rect 41337 2397 41371 2431
rect 43269 2397 43303 2431
rect 45845 2397 45879 2431
rect 47777 2397 47811 2431
rect 22845 2329 22879 2363
rect 25053 2329 25087 2363
rect 28549 2329 28583 2363
rect 29837 2261 29871 2295
<< metal1 >>
rect 19702 47744 19708 47796
rect 19760 47784 19766 47796
rect 22370 47784 22376 47796
rect 19760 47756 22376 47784
rect 19760 47744 19766 47756
rect 22370 47744 22376 47756
rect 22428 47744 22434 47796
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 4706 47240 4712 47252
rect 4667 47212 4712 47240
rect 4706 47200 4712 47212
rect 4764 47200 4770 47252
rect 5353 47243 5411 47249
rect 5353 47209 5365 47243
rect 5399 47240 5411 47243
rect 5810 47240 5816 47252
rect 5399 47212 5816 47240
rect 5399 47209 5411 47212
rect 5353 47203 5411 47209
rect 5810 47200 5816 47212
rect 5868 47200 5874 47252
rect 5994 47240 6000 47252
rect 5955 47212 6000 47240
rect 5994 47200 6000 47212
rect 6052 47200 6058 47252
rect 7098 47240 7104 47252
rect 7059 47212 7104 47240
rect 7098 47200 7104 47212
rect 7156 47200 7162 47252
rect 7742 47240 7748 47252
rect 7703 47212 7748 47240
rect 7742 47200 7748 47212
rect 7800 47200 7806 47252
rect 8386 47240 8392 47252
rect 8347 47212 8392 47240
rect 8386 47200 8392 47212
rect 8444 47200 8450 47252
rect 9122 47240 9128 47252
rect 9083 47212 9128 47240
rect 9122 47200 9128 47212
rect 9180 47200 9186 47252
rect 10226 47240 10232 47252
rect 10187 47212 10232 47240
rect 10226 47200 10232 47212
rect 10284 47200 10290 47252
rect 11146 47240 11152 47252
rect 11107 47212 11152 47240
rect 11146 47200 11152 47212
rect 11204 47200 11210 47252
rect 12434 47200 12440 47252
rect 12492 47240 12498 47252
rect 13538 47240 13544 47252
rect 12492 47212 12537 47240
rect 13499 47212 13544 47240
rect 12492 47200 12498 47212
rect 13538 47200 13544 47212
rect 13596 47200 13602 47252
rect 15013 47243 15071 47249
rect 15013 47209 15025 47243
rect 15059 47240 15071 47243
rect 16850 47240 16856 47252
rect 15059 47212 16856 47240
rect 15059 47209 15071 47212
rect 15013 47203 15071 47209
rect 16850 47200 16856 47212
rect 16908 47200 16914 47252
rect 20162 47240 20168 47252
rect 17236 47212 20168 47240
rect 15657 47107 15715 47113
rect 15657 47073 15669 47107
rect 15703 47104 15715 47107
rect 17236 47104 17264 47212
rect 20162 47200 20168 47212
rect 20220 47200 20226 47252
rect 20622 47240 20628 47252
rect 20583 47212 20628 47240
rect 20622 47200 20628 47212
rect 20680 47200 20686 47252
rect 24029 47243 24087 47249
rect 24029 47209 24041 47243
rect 24075 47240 24087 47243
rect 25682 47240 25688 47252
rect 24075 47212 25688 47240
rect 24075 47209 24087 47212
rect 24029 47203 24087 47209
rect 25682 47200 25688 47212
rect 25740 47200 25746 47252
rect 26050 47240 26056 47252
rect 26011 47212 26056 47240
rect 26050 47200 26056 47212
rect 26108 47200 26114 47252
rect 40402 47200 40408 47252
rect 40460 47240 40466 47252
rect 43901 47243 43959 47249
rect 43901 47240 43913 47243
rect 40460 47212 43913 47240
rect 40460 47200 40466 47212
rect 43901 47209 43913 47212
rect 43947 47209 43959 47243
rect 43901 47203 43959 47209
rect 44174 47200 44180 47252
rect 44232 47240 44238 47252
rect 45189 47243 45247 47249
rect 45189 47240 45201 47243
rect 44232 47212 45201 47240
rect 44232 47200 44238 47212
rect 45189 47209 45201 47212
rect 45235 47209 45247 47243
rect 45189 47203 45247 47209
rect 45922 47200 45928 47252
rect 45980 47240 45986 47252
rect 46477 47243 46535 47249
rect 46477 47240 46489 47243
rect 45980 47212 46489 47240
rect 45980 47200 45986 47212
rect 46477 47209 46489 47212
rect 46523 47209 46535 47243
rect 46477 47203 46535 47209
rect 19702 47172 19708 47184
rect 15703 47076 17264 47104
rect 17420 47144 19708 47172
rect 15703 47073 15715 47076
rect 15657 47067 15715 47073
rect 16301 47039 16359 47045
rect 16301 47005 16313 47039
rect 16347 47036 16359 47039
rect 17420 47036 17448 47144
rect 19702 47132 19708 47144
rect 19760 47132 19766 47184
rect 19886 47132 19892 47184
rect 19944 47172 19950 47184
rect 33870 47172 33876 47184
rect 19944 47144 24624 47172
rect 19944 47132 19950 47144
rect 24596 47113 24624 47144
rect 33244 47144 33876 47172
rect 19429 47107 19487 47113
rect 19429 47104 19441 47107
rect 17512 47076 19441 47104
rect 17512 47045 17540 47076
rect 19429 47073 19441 47076
rect 19475 47073 19487 47107
rect 19429 47067 19487 47073
rect 19981 47107 20039 47113
rect 19981 47073 19993 47107
rect 20027 47073 20039 47107
rect 22557 47107 22615 47113
rect 22557 47104 22569 47107
rect 19981 47067 20039 47073
rect 21744 47076 22569 47104
rect 16347 47008 17448 47036
rect 17497 47039 17555 47045
rect 16347 47005 16359 47008
rect 16301 46999 16359 47005
rect 17497 47005 17509 47039
rect 17543 47005 17555 47039
rect 17497 46999 17555 47005
rect 18417 47039 18475 47045
rect 18417 47005 18429 47039
rect 18463 47005 18475 47039
rect 18417 46999 18475 47005
rect 18509 47039 18567 47045
rect 18509 47005 18521 47039
rect 18555 47036 18567 47039
rect 18690 47036 18696 47048
rect 18555 47008 18696 47036
rect 18555 47005 18567 47008
rect 18509 46999 18567 47005
rect 17957 46971 18015 46977
rect 17328 46940 17908 46968
rect 10594 46860 10600 46912
rect 10652 46900 10658 46912
rect 17126 46900 17132 46912
rect 10652 46872 17132 46900
rect 10652 46860 10658 46872
rect 17126 46860 17132 46872
rect 17184 46860 17190 46912
rect 17328 46909 17356 46940
rect 17313 46903 17371 46909
rect 17313 46869 17325 46903
rect 17359 46869 17371 46903
rect 17880 46900 17908 46940
rect 17957 46937 17969 46971
rect 18003 46968 18015 46971
rect 18138 46968 18144 46980
rect 18003 46940 18144 46968
rect 18003 46937 18015 46940
rect 17957 46931 18015 46937
rect 18138 46928 18144 46940
rect 18196 46928 18202 46980
rect 18432 46968 18460 46999
rect 18690 46996 18696 47008
rect 18748 47036 18754 47048
rect 19886 47036 19892 47048
rect 18748 47008 19334 47036
rect 19847 47008 19892 47036
rect 18748 46996 18754 47008
rect 18966 46968 18972 46980
rect 18432 46940 18972 46968
rect 18966 46928 18972 46940
rect 19024 46928 19030 46980
rect 19306 46968 19334 47008
rect 19886 46996 19892 47008
rect 19944 46996 19950 47048
rect 19996 46968 20024 47067
rect 20438 47036 20444 47048
rect 20399 47008 20444 47036
rect 20438 46996 20444 47008
rect 20496 46996 20502 47048
rect 21453 47039 21511 47045
rect 21453 47005 21465 47039
rect 21499 47036 21511 47039
rect 21744 47036 21772 47076
rect 22557 47073 22569 47076
rect 22603 47073 22615 47107
rect 22557 47067 22615 47073
rect 24581 47107 24639 47113
rect 24581 47073 24593 47107
rect 24627 47073 24639 47107
rect 27798 47104 27804 47116
rect 24581 47067 24639 47073
rect 25424 47076 27804 47104
rect 21499 47008 21772 47036
rect 22005 47039 22063 47045
rect 21499 47005 21511 47008
rect 21453 46999 21511 47005
rect 22005 47005 22017 47039
rect 22051 47005 22063 47039
rect 22005 46999 22063 47005
rect 22020 46968 22048 46999
rect 22094 46996 22100 47048
rect 22152 47036 22158 47048
rect 23385 47039 23443 47045
rect 22152 47008 22197 47036
rect 22152 46996 22158 47008
rect 23385 47005 23397 47039
rect 23431 47005 23443 47039
rect 25130 47036 25136 47048
rect 25091 47008 25136 47036
rect 23385 46999 23443 47005
rect 19306 46940 22048 46968
rect 23400 46968 23428 46999
rect 25130 46996 25136 47008
rect 25188 46996 25194 47048
rect 25424 47045 25452 47076
rect 27798 47064 27804 47076
rect 27856 47064 27862 47116
rect 29733 47107 29791 47113
rect 29733 47104 29745 47107
rect 28000 47076 29745 47104
rect 25409 47039 25467 47045
rect 25409 47005 25421 47039
rect 25455 47005 25467 47039
rect 25590 47036 25596 47048
rect 25551 47008 25596 47036
rect 25409 46999 25467 47005
rect 25590 46996 25596 47008
rect 25648 46996 25654 47048
rect 27706 47036 27712 47048
rect 27667 47008 27712 47036
rect 27706 46996 27712 47008
rect 27764 46996 27770 47048
rect 28000 47045 28028 47076
rect 29733 47073 29745 47076
rect 29779 47104 29791 47107
rect 30282 47104 30288 47116
rect 29779 47076 30288 47104
rect 29779 47073 29791 47076
rect 29733 47067 29791 47073
rect 30282 47064 30288 47076
rect 30340 47064 30346 47116
rect 31202 47104 31208 47116
rect 31163 47076 31208 47104
rect 31202 47064 31208 47076
rect 31260 47064 31266 47116
rect 33244 47113 33272 47144
rect 33870 47132 33876 47144
rect 33928 47172 33934 47184
rect 36354 47172 36360 47184
rect 33928 47144 36360 47172
rect 33928 47132 33934 47144
rect 36354 47132 36360 47144
rect 36412 47172 36418 47184
rect 36814 47172 36820 47184
rect 36412 47144 36820 47172
rect 36412 47132 36418 47144
rect 36814 47132 36820 47144
rect 36872 47132 36878 47184
rect 38197 47175 38255 47181
rect 38197 47141 38209 47175
rect 38243 47141 38255 47175
rect 38197 47135 38255 47141
rect 33229 47107 33287 47113
rect 33229 47073 33241 47107
rect 33275 47073 33287 47107
rect 37642 47104 37648 47116
rect 33229 47067 33287 47073
rect 33520 47076 37648 47104
rect 27985 47039 28043 47045
rect 27985 47005 27997 47039
rect 28031 47005 28043 47039
rect 27985 46999 28043 47005
rect 28169 47039 28227 47045
rect 28169 47005 28181 47039
rect 28215 47005 28227 47039
rect 28902 47036 28908 47048
rect 28863 47008 28908 47036
rect 28169 46999 28227 47005
rect 26878 46968 26884 46980
rect 23400 46940 26884 46968
rect 21468 46912 21496 46940
rect 26878 46928 26884 46940
rect 26936 46928 26942 46980
rect 27154 46968 27160 46980
rect 27115 46940 27160 46968
rect 27154 46928 27160 46940
rect 27212 46928 27218 46980
rect 18414 46900 18420 46912
rect 17880 46872 18420 46900
rect 17313 46863 17371 46869
rect 18414 46860 18420 46872
rect 18472 46860 18478 46912
rect 18598 46860 18604 46912
rect 18656 46900 18662 46912
rect 21174 46900 21180 46912
rect 18656 46872 21180 46900
rect 18656 46860 18662 46872
rect 21174 46860 21180 46872
rect 21232 46900 21238 46912
rect 21269 46903 21327 46909
rect 21269 46900 21281 46903
rect 21232 46872 21281 46900
rect 21232 46860 21238 46872
rect 21269 46869 21281 46872
rect 21315 46869 21327 46903
rect 21269 46863 21327 46869
rect 21450 46860 21456 46912
rect 21508 46860 21514 46912
rect 24210 46860 24216 46912
rect 24268 46900 24274 46912
rect 26418 46900 26424 46912
rect 24268 46872 26424 46900
rect 24268 46860 24274 46872
rect 26418 46860 26424 46872
rect 26476 46900 26482 46912
rect 28000 46900 28028 46999
rect 28184 46968 28212 46999
rect 28902 46996 28908 47008
rect 28960 47036 28966 47048
rect 30006 47036 30012 47048
rect 28960 47008 30012 47036
rect 28960 46996 28966 47008
rect 30006 46996 30012 47008
rect 30064 46996 30070 47048
rect 30745 47039 30803 47045
rect 30745 47005 30757 47039
rect 30791 47036 30803 47039
rect 30834 47036 30840 47048
rect 30791 47008 30840 47036
rect 30791 47005 30803 47008
rect 30745 46999 30803 47005
rect 30834 46996 30840 47008
rect 30892 46996 30898 47048
rect 31113 47039 31171 47045
rect 31113 47005 31125 47039
rect 31159 47036 31171 47039
rect 31294 47036 31300 47048
rect 31159 47008 31300 47036
rect 31159 47005 31171 47008
rect 31113 46999 31171 47005
rect 31294 46996 31300 47008
rect 31352 46996 31358 47048
rect 33520 47045 33548 47076
rect 33505 47039 33563 47045
rect 33505 47005 33517 47039
rect 33551 47005 33563 47039
rect 33686 47036 33692 47048
rect 33647 47008 33692 47036
rect 33505 46999 33563 47005
rect 30285 46971 30343 46977
rect 28184 46940 29132 46968
rect 29104 46909 29132 46940
rect 30285 46937 30297 46971
rect 30331 46968 30343 46971
rect 30374 46968 30380 46980
rect 30331 46940 30380 46968
rect 30331 46937 30343 46940
rect 30285 46931 30343 46937
rect 30374 46928 30380 46940
rect 30432 46928 30438 46980
rect 32030 46928 32036 46980
rect 32088 46968 32094 46980
rect 32677 46971 32735 46977
rect 32677 46968 32689 46971
rect 32088 46940 32689 46968
rect 32088 46928 32094 46940
rect 32677 46937 32689 46940
rect 32723 46937 32735 46971
rect 32677 46931 32735 46937
rect 33134 46928 33140 46980
rect 33192 46968 33198 46980
rect 33520 46968 33548 46999
rect 33686 46996 33692 47008
rect 33744 46996 33750 47048
rect 34149 47039 34207 47045
rect 34149 47005 34161 47039
rect 34195 47005 34207 47039
rect 34149 46999 34207 47005
rect 35345 47039 35403 47045
rect 35345 47005 35357 47039
rect 35391 47005 35403 47039
rect 35526 47036 35532 47048
rect 35487 47008 35532 47036
rect 35345 46999 35403 47005
rect 33192 46940 33548 46968
rect 33192 46928 33198 46940
rect 26476 46872 28028 46900
rect 29089 46903 29147 46909
rect 26476 46860 26482 46872
rect 29089 46869 29101 46903
rect 29135 46900 29147 46903
rect 29362 46900 29368 46912
rect 29135 46872 29368 46900
rect 29135 46869 29147 46872
rect 29089 46863 29147 46869
rect 29362 46860 29368 46872
rect 29420 46860 29426 46912
rect 29822 46860 29828 46912
rect 29880 46900 29886 46912
rect 34164 46900 34192 46999
rect 34422 46928 34428 46980
rect 34480 46968 34486 46980
rect 34885 46971 34943 46977
rect 34885 46968 34897 46971
rect 34480 46940 34897 46968
rect 34480 46928 34486 46940
rect 34885 46937 34897 46940
rect 34931 46937 34943 46971
rect 35360 46968 35388 46999
rect 35526 46996 35532 47008
rect 35584 46996 35590 47048
rect 35728 47045 35756 47076
rect 37642 47064 37648 47076
rect 37700 47104 37706 47116
rect 38212 47104 38240 47135
rect 38470 47132 38476 47184
rect 38528 47172 38534 47184
rect 38933 47175 38991 47181
rect 38933 47172 38945 47175
rect 38528 47144 38945 47172
rect 38528 47132 38534 47144
rect 38933 47141 38945 47144
rect 38979 47141 38991 47175
rect 38933 47135 38991 47141
rect 41417 47175 41475 47181
rect 41417 47141 41429 47175
rect 41463 47172 41475 47175
rect 41782 47172 41788 47184
rect 41463 47144 41788 47172
rect 41463 47141 41475 47144
rect 41417 47135 41475 47141
rect 41782 47132 41788 47144
rect 41840 47132 41846 47184
rect 44266 47132 44272 47184
rect 44324 47172 44330 47184
rect 44545 47175 44603 47181
rect 44545 47172 44557 47175
rect 44324 47144 44557 47172
rect 44324 47132 44330 47144
rect 44545 47141 44557 47144
rect 44591 47141 44603 47175
rect 44545 47135 44603 47141
rect 37700 47076 38240 47104
rect 37700 47064 37706 47076
rect 35713 47039 35771 47045
rect 35713 47005 35725 47039
rect 35759 47005 35771 47039
rect 36354 47036 36360 47048
rect 36315 47008 36360 47036
rect 35713 46999 35771 47005
rect 36354 46996 36360 47008
rect 36412 46996 36418 47048
rect 37458 47036 37464 47048
rect 37419 47008 37464 47036
rect 37458 46996 37464 47008
rect 37516 46996 37522 47048
rect 38378 47036 38384 47048
rect 38339 47008 38384 47036
rect 38378 46996 38384 47008
rect 38436 46996 38442 47048
rect 38654 46996 38660 47048
rect 38712 47036 38718 47048
rect 39117 47039 39175 47045
rect 39117 47036 39129 47039
rect 38712 47008 39129 47036
rect 38712 46996 38718 47008
rect 39117 47005 39129 47008
rect 39163 47005 39175 47039
rect 39117 46999 39175 47005
rect 40218 46996 40224 47048
rect 40276 47036 40282 47048
rect 40865 47039 40923 47045
rect 40865 47036 40877 47039
rect 40276 47008 40877 47036
rect 40276 46996 40282 47008
rect 40865 47005 40877 47008
rect 40911 47036 40923 47039
rect 41601 47039 41659 47045
rect 41601 47036 41613 47039
rect 40911 47008 41613 47036
rect 40911 47005 40923 47008
rect 40865 46999 40923 47005
rect 41601 47005 41613 47008
rect 41647 47005 41659 47039
rect 41601 46999 41659 47005
rect 36630 46968 36636 46980
rect 35360 46940 36636 46968
rect 34885 46931 34943 46937
rect 36630 46928 36636 46940
rect 36688 46968 36694 46980
rect 39390 46968 39396 46980
rect 36688 46940 37228 46968
rect 36688 46928 36694 46940
rect 29880 46872 34192 46900
rect 29880 46860 29886 46872
rect 35526 46860 35532 46912
rect 35584 46900 35590 46912
rect 35710 46900 35716 46912
rect 35584 46872 35716 46900
rect 35584 46860 35590 46872
rect 35710 46860 35716 46872
rect 35768 46860 35774 46912
rect 35986 46860 35992 46912
rect 36044 46900 36050 46912
rect 37090 46900 37096 46912
rect 36044 46872 37096 46900
rect 36044 46860 36050 46872
rect 37090 46860 37096 46872
rect 37148 46860 37154 46912
rect 37200 46900 37228 46940
rect 37752 46940 39396 46968
rect 37752 46900 37780 46940
rect 39390 46928 39396 46940
rect 39448 46928 39454 46980
rect 37200 46872 37780 46900
rect 37826 46860 37832 46912
rect 37884 46900 37890 46912
rect 39942 46900 39948 46912
rect 37884 46872 39948 46900
rect 37884 46860 37890 46872
rect 39942 46860 39948 46872
rect 40000 46860 40006 46912
rect 40586 46900 40592 46912
rect 40547 46872 40592 46900
rect 40586 46860 40592 46872
rect 40644 46860 40650 46912
rect 41616 46900 41644 46999
rect 42426 46996 42432 47048
rect 42484 47036 42490 47048
rect 42613 47039 42671 47045
rect 42613 47036 42625 47039
rect 42484 47008 42625 47036
rect 42484 46996 42490 47008
rect 42613 47005 42625 47008
rect 42659 47005 42671 47039
rect 43254 47036 43260 47048
rect 43215 47008 43260 47036
rect 42613 46999 42671 47005
rect 43254 46996 43260 47008
rect 43312 46996 43318 47048
rect 45833 47039 45891 47045
rect 45833 47036 45845 47039
rect 45526 47008 45845 47036
rect 43898 46900 43904 46912
rect 41616 46872 43904 46900
rect 43898 46860 43904 46872
rect 43956 46860 43962 46912
rect 44726 46860 44732 46912
rect 44784 46900 44790 46912
rect 45526 46900 45554 47008
rect 45833 47005 45845 47008
rect 45879 47005 45891 47039
rect 45833 46999 45891 47005
rect 44784 46872 45554 46900
rect 44784 46860 44790 46872
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 16114 46696 16120 46708
rect 16075 46668 16120 46696
rect 16114 46656 16120 46668
rect 16172 46656 16178 46708
rect 17218 46656 17224 46708
rect 17276 46656 17282 46708
rect 21634 46696 21640 46708
rect 18800 46668 21640 46696
rect 9490 46588 9496 46640
rect 9548 46628 9554 46640
rect 17236 46628 17264 46656
rect 9548 46600 12434 46628
rect 17236 46600 18276 46628
rect 9548 46588 9554 46600
rect 6914 46520 6920 46572
rect 6972 46560 6978 46572
rect 6972 46532 7017 46560
rect 6972 46520 6978 46532
rect 12406 46356 12434 46600
rect 14642 46560 14648 46572
rect 14603 46532 14648 46560
rect 14642 46520 14648 46532
rect 14700 46520 14706 46572
rect 15562 46560 15568 46572
rect 15523 46532 15568 46560
rect 15562 46520 15568 46532
rect 15620 46520 15626 46572
rect 16301 46563 16359 46569
rect 16301 46529 16313 46563
rect 16347 46560 16359 46563
rect 17221 46563 17279 46569
rect 17221 46560 17233 46563
rect 16347 46532 17233 46560
rect 16347 46529 16359 46532
rect 16301 46523 16359 46529
rect 17221 46529 17233 46532
rect 17267 46529 17279 46563
rect 17221 46523 17279 46529
rect 17402 46520 17408 46572
rect 17460 46560 17466 46572
rect 17681 46563 17739 46569
rect 17681 46560 17693 46563
rect 17460 46532 17693 46560
rect 17460 46520 17466 46532
rect 17681 46529 17693 46532
rect 17727 46560 17739 46563
rect 18046 46560 18052 46572
rect 17727 46532 18052 46560
rect 17727 46529 17739 46532
rect 17681 46523 17739 46529
rect 18046 46520 18052 46532
rect 18104 46520 18110 46572
rect 18248 46569 18276 46600
rect 18233 46563 18291 46569
rect 18233 46529 18245 46563
rect 18279 46560 18291 46563
rect 18322 46560 18328 46572
rect 18279 46532 18328 46560
rect 18279 46529 18291 46532
rect 18233 46523 18291 46529
rect 18322 46520 18328 46532
rect 18380 46520 18386 46572
rect 18414 46520 18420 46572
rect 18472 46560 18478 46572
rect 18800 46560 18828 46668
rect 21634 46656 21640 46668
rect 21692 46656 21698 46708
rect 30374 46696 30380 46708
rect 24136 46668 30380 46696
rect 19978 46628 19984 46640
rect 19168 46600 19984 46628
rect 18966 46560 18972 46572
rect 18472 46532 18828 46560
rect 18927 46532 18972 46560
rect 18472 46520 18478 46532
rect 18966 46520 18972 46532
rect 19024 46520 19030 46572
rect 19168 46569 19196 46600
rect 19978 46588 19984 46600
rect 20036 46588 20042 46640
rect 21726 46628 21732 46640
rect 21376 46600 21732 46628
rect 19153 46563 19211 46569
rect 19153 46529 19165 46563
rect 19199 46529 19211 46563
rect 19153 46523 19211 46529
rect 19886 46520 19892 46572
rect 19944 46560 19950 46572
rect 20165 46563 20223 46569
rect 20165 46560 20177 46563
rect 19944 46532 20177 46560
rect 19944 46520 19950 46532
rect 20165 46529 20177 46532
rect 20211 46560 20223 46563
rect 20438 46560 20444 46572
rect 20211 46532 20444 46560
rect 20211 46529 20223 46532
rect 20165 46523 20223 46529
rect 20438 46520 20444 46532
rect 20496 46520 20502 46572
rect 21376 46569 21404 46600
rect 21726 46588 21732 46600
rect 21784 46588 21790 46640
rect 23842 46628 23848 46640
rect 23584 46600 23848 46628
rect 21361 46563 21419 46569
rect 21361 46529 21373 46563
rect 21407 46529 21419 46563
rect 21361 46523 21419 46529
rect 22094 46520 22100 46572
rect 22152 46560 22158 46572
rect 22830 46560 22836 46572
rect 22152 46532 22197 46560
rect 22791 46532 22836 46560
rect 22152 46520 22158 46532
rect 22830 46520 22836 46532
rect 22888 46520 22894 46572
rect 23468 46563 23526 46569
rect 23468 46529 23480 46563
rect 23514 46560 23526 46563
rect 23584 46560 23612 46600
rect 23842 46588 23848 46600
rect 23900 46588 23906 46640
rect 24136 46628 24164 46668
rect 30374 46656 30380 46668
rect 30432 46656 30438 46708
rect 32674 46656 32680 46708
rect 32732 46696 32738 46708
rect 34146 46696 34152 46708
rect 32732 46668 34152 46696
rect 32732 46656 32738 46668
rect 34146 46656 34152 46668
rect 34204 46656 34210 46708
rect 37458 46696 37464 46708
rect 34256 46668 37464 46696
rect 24044 46600 24164 46628
rect 25869 46631 25927 46637
rect 24044 46569 24072 46600
rect 25869 46597 25881 46631
rect 25915 46628 25927 46631
rect 27154 46628 27160 46640
rect 25915 46600 27160 46628
rect 25915 46597 25927 46600
rect 25869 46591 25927 46597
rect 27154 46588 27160 46600
rect 27212 46588 27218 46640
rect 27798 46628 27804 46640
rect 27759 46600 27804 46628
rect 27798 46588 27804 46600
rect 27856 46588 27862 46640
rect 28920 46600 30512 46628
rect 23514 46532 23612 46560
rect 23661 46563 23719 46569
rect 23514 46529 23526 46532
rect 23468 46523 23526 46529
rect 23661 46529 23673 46563
rect 23707 46529 23719 46563
rect 23661 46523 23719 46529
rect 24029 46563 24087 46569
rect 24029 46529 24041 46563
rect 24075 46529 24087 46563
rect 24029 46523 24087 46529
rect 13906 46452 13912 46504
rect 13964 46492 13970 46504
rect 17586 46492 17592 46504
rect 13964 46464 17592 46492
rect 13964 46452 13970 46464
rect 17586 46452 17592 46464
rect 17644 46452 17650 46504
rect 17773 46495 17831 46501
rect 17773 46461 17785 46495
rect 17819 46492 17831 46495
rect 18598 46492 18604 46504
rect 17819 46464 18604 46492
rect 17819 46461 17831 46464
rect 17773 46455 17831 46461
rect 18598 46452 18604 46464
rect 18656 46452 18662 46504
rect 19426 46452 19432 46504
rect 19484 46452 19490 46504
rect 20898 46492 20904 46504
rect 20859 46464 20904 46492
rect 20898 46452 20904 46464
rect 20956 46452 20962 46504
rect 21450 46452 21456 46504
rect 21508 46501 21514 46504
rect 21508 46492 21515 46501
rect 23676 46492 23704 46523
rect 24118 46520 24124 46572
rect 24176 46560 24182 46572
rect 24302 46560 24308 46572
rect 24176 46532 24221 46560
rect 24263 46532 24308 46560
rect 24176 46520 24182 46532
rect 24302 46520 24308 46532
rect 24360 46520 24366 46572
rect 25590 46520 25596 46572
rect 25648 46560 25654 46572
rect 26237 46563 26295 46569
rect 26237 46560 26249 46563
rect 25648 46532 26249 46560
rect 25648 46520 25654 46532
rect 26237 46529 26249 46532
rect 26283 46529 26295 46563
rect 26237 46523 26295 46529
rect 26329 46563 26387 46569
rect 26329 46529 26341 46563
rect 26375 46560 26387 46563
rect 26970 46560 26976 46572
rect 26375 46532 26976 46560
rect 26375 46529 26387 46532
rect 26329 46523 26387 46529
rect 26970 46520 26976 46532
rect 27028 46520 27034 46572
rect 27062 46520 27068 46572
rect 27120 46560 27126 46572
rect 28920 46560 28948 46600
rect 30484 46572 30512 46600
rect 31570 46588 31576 46640
rect 31628 46628 31634 46640
rect 33502 46628 33508 46640
rect 31628 46600 33508 46628
rect 31628 46588 31634 46600
rect 33502 46588 33508 46600
rect 33560 46588 33566 46640
rect 33594 46588 33600 46640
rect 33652 46628 33658 46640
rect 33689 46631 33747 46637
rect 33689 46628 33701 46631
rect 33652 46600 33701 46628
rect 33652 46588 33658 46600
rect 33689 46597 33701 46600
rect 33735 46597 33747 46631
rect 33689 46591 33747 46597
rect 29086 46560 29092 46572
rect 27120 46532 28948 46560
rect 29047 46532 29092 46560
rect 27120 46520 27126 46532
rect 29086 46520 29092 46532
rect 29144 46520 29150 46572
rect 29638 46560 29644 46572
rect 29599 46532 29644 46560
rect 29638 46520 29644 46532
rect 29696 46520 29702 46572
rect 30466 46560 30472 46572
rect 30379 46532 30472 46560
rect 30466 46520 30472 46532
rect 30524 46520 30530 46572
rect 31294 46560 31300 46572
rect 31255 46532 31300 46560
rect 31294 46520 31300 46532
rect 31352 46520 31358 46572
rect 33045 46563 33103 46569
rect 33045 46529 33057 46563
rect 33091 46560 33103 46563
rect 33134 46560 33140 46572
rect 33091 46532 33140 46560
rect 33091 46529 33103 46532
rect 33045 46523 33103 46529
rect 33134 46520 33140 46532
rect 33192 46520 33198 46572
rect 33226 46520 33232 46572
rect 33284 46560 33290 46572
rect 34149 46563 34207 46569
rect 34149 46560 34161 46563
rect 33284 46532 33329 46560
rect 33520 46532 34161 46560
rect 33284 46520 33290 46532
rect 30932 46504 30984 46510
rect 26418 46492 26424 46504
rect 21508 46464 21553 46492
rect 22204 46464 25544 46492
rect 26379 46464 26424 46492
rect 21508 46455 21515 46464
rect 21508 46452 21514 46455
rect 15010 46384 15016 46436
rect 15068 46424 15074 46436
rect 19334 46424 19340 46436
rect 15068 46396 19340 46424
rect 15068 46384 15074 46396
rect 19334 46384 19340 46396
rect 19392 46384 19398 46436
rect 19444 46424 19472 46452
rect 22204 46424 22232 46464
rect 19444 46396 22232 46424
rect 22281 46427 22339 46433
rect 22281 46393 22293 46427
rect 22327 46424 22339 46427
rect 22738 46424 22744 46436
rect 22327 46396 22744 46424
rect 22327 46393 22339 46396
rect 22281 46387 22339 46393
rect 22738 46384 22744 46396
rect 22796 46384 22802 46436
rect 25406 46424 25412 46436
rect 25367 46396 25412 46424
rect 25406 46384 25412 46396
rect 25464 46384 25470 46436
rect 25516 46424 25544 46464
rect 26418 46452 26424 46464
rect 26476 46452 26482 46504
rect 26786 46452 26792 46504
rect 26844 46492 26850 46504
rect 27157 46495 27215 46501
rect 27157 46492 27169 46495
rect 26844 46464 27169 46492
rect 26844 46452 26850 46464
rect 27157 46461 27169 46464
rect 27203 46461 27215 46495
rect 27157 46455 27215 46461
rect 31110 46492 31116 46504
rect 31071 46464 31116 46492
rect 31110 46452 31116 46464
rect 31168 46452 31174 46504
rect 32769 46495 32827 46501
rect 32769 46461 32781 46495
rect 32815 46492 32827 46495
rect 33520 46492 33548 46532
rect 34149 46529 34161 46532
rect 34195 46529 34207 46563
rect 34149 46523 34207 46529
rect 32815 46464 33548 46492
rect 32815 46461 32827 46464
rect 32769 46455 32827 46461
rect 30932 46446 30984 46452
rect 30285 46427 30343 46433
rect 30285 46424 30297 46427
rect 25516 46396 30297 46424
rect 30285 46393 30297 46396
rect 30331 46393 30343 46427
rect 30285 46387 30343 46393
rect 32306 46384 32312 46436
rect 32364 46424 32370 46436
rect 34256 46424 34284 46668
rect 37458 46656 37464 46668
rect 37516 46656 37522 46708
rect 38194 46656 38200 46708
rect 38252 46696 38258 46708
rect 41414 46696 41420 46708
rect 38252 46668 41420 46696
rect 38252 46656 38258 46668
rect 41414 46656 41420 46668
rect 41472 46656 41478 46708
rect 34624 46600 36676 46628
rect 34624 46572 34652 46600
rect 34422 46560 34428 46572
rect 34383 46532 34428 46560
rect 34422 46520 34428 46532
rect 34480 46520 34486 46572
rect 34606 46560 34612 46572
rect 34567 46532 34612 46560
rect 34606 46520 34612 46532
rect 34664 46520 34670 46572
rect 35161 46563 35219 46569
rect 35161 46529 35173 46563
rect 35207 46560 35219 46563
rect 35342 46560 35348 46572
rect 35207 46532 35348 46560
rect 35207 46529 35219 46532
rect 35161 46523 35219 46529
rect 35342 46520 35348 46532
rect 35400 46520 35406 46572
rect 35526 46520 35532 46572
rect 35584 46560 35590 46572
rect 35621 46563 35679 46569
rect 35621 46560 35633 46563
rect 35584 46532 35633 46560
rect 35584 46520 35590 46532
rect 35621 46529 35633 46532
rect 35667 46529 35679 46563
rect 35621 46523 35679 46529
rect 36449 46563 36507 46569
rect 36449 46529 36461 46563
rect 36495 46529 36507 46563
rect 36449 46523 36507 46529
rect 34790 46492 34796 46504
rect 34751 46464 34796 46492
rect 34790 46452 34796 46464
rect 34848 46452 34854 46504
rect 36173 46495 36231 46501
rect 36173 46461 36185 46495
rect 36219 46492 36231 46495
rect 36354 46492 36360 46504
rect 36219 46464 36360 46492
rect 36219 46461 36231 46464
rect 36173 46455 36231 46461
rect 36354 46452 36360 46464
rect 36412 46452 36418 46504
rect 36262 46424 36268 46436
rect 32364 46396 34284 46424
rect 34440 46396 36268 46424
rect 32364 46384 32370 46396
rect 18782 46356 18788 46368
rect 12406 46328 18788 46356
rect 18782 46316 18788 46328
rect 18840 46316 18846 46368
rect 19426 46356 19432 46368
rect 19387 46328 19432 46356
rect 19426 46316 19432 46328
rect 19484 46316 19490 46368
rect 19978 46316 19984 46368
rect 20036 46356 20042 46368
rect 20349 46359 20407 46365
rect 20349 46356 20361 46359
rect 20036 46328 20361 46356
rect 20036 46316 20042 46328
rect 20349 46325 20361 46328
rect 20395 46356 20407 46359
rect 24854 46356 24860 46368
rect 20395 46328 24860 46356
rect 20395 46325 20407 46328
rect 20349 46319 20407 46325
rect 24854 46316 24860 46328
rect 24912 46316 24918 46368
rect 24949 46359 25007 46365
rect 24949 46325 24961 46359
rect 24995 46356 25007 46359
rect 26234 46356 26240 46368
rect 24995 46328 26240 46356
rect 24995 46325 25007 46328
rect 24949 46319 25007 46325
rect 26234 46316 26240 46328
rect 26292 46316 26298 46368
rect 33042 46316 33048 46368
rect 33100 46356 33106 46368
rect 34440 46356 34468 46396
rect 36262 46384 36268 46396
rect 36320 46384 36326 46436
rect 36464 46424 36492 46523
rect 36648 46504 36676 46600
rect 36814 46588 36820 46640
rect 36872 46628 36878 46640
rect 41969 46631 42027 46637
rect 41969 46628 41981 46631
rect 36872 46600 41981 46628
rect 36872 46588 36878 46600
rect 41969 46597 41981 46600
rect 42015 46597 42027 46631
rect 41969 46591 42027 46597
rect 38289 46563 38347 46569
rect 38289 46529 38301 46563
rect 38335 46529 38347 46563
rect 38470 46560 38476 46572
rect 38431 46532 38476 46560
rect 38289 46523 38347 46529
rect 36630 46492 36636 46504
rect 36591 46464 36636 46492
rect 36630 46452 36636 46464
rect 36688 46452 36694 46504
rect 36906 46452 36912 46504
rect 36964 46492 36970 46504
rect 37461 46495 37519 46501
rect 37461 46492 37473 46495
rect 36964 46464 37473 46492
rect 36964 46452 36970 46464
rect 37461 46461 37473 46464
rect 37507 46461 37519 46495
rect 37461 46455 37519 46461
rect 38013 46495 38071 46501
rect 38013 46461 38025 46495
rect 38059 46492 38071 46495
rect 38102 46492 38108 46504
rect 38059 46464 38108 46492
rect 38059 46461 38071 46464
rect 38013 46455 38071 46461
rect 38102 46452 38108 46464
rect 38160 46452 38166 46504
rect 38304 46492 38332 46523
rect 38470 46520 38476 46532
rect 38528 46520 38534 46572
rect 39574 46560 39580 46572
rect 38672 46532 39580 46560
rect 38378 46492 38384 46504
rect 38291 46464 38384 46492
rect 38378 46452 38384 46464
rect 38436 46492 38442 46504
rect 38672 46492 38700 46532
rect 39574 46520 39580 46532
rect 39632 46520 39638 46572
rect 40218 46560 40224 46572
rect 40179 46532 40224 46560
rect 40218 46520 40224 46532
rect 40276 46520 40282 46572
rect 40310 46520 40316 46572
rect 40368 46560 40374 46572
rect 43257 46563 43315 46569
rect 43257 46560 43269 46563
rect 40368 46532 43269 46560
rect 40368 46520 40374 46532
rect 43257 46529 43269 46532
rect 43303 46529 43315 46563
rect 43257 46523 43315 46529
rect 43346 46520 43352 46572
rect 43404 46560 43410 46572
rect 44545 46563 44603 46569
rect 44545 46560 44557 46563
rect 43404 46532 44557 46560
rect 43404 46520 43410 46532
rect 44545 46529 44557 46532
rect 44591 46529 44603 46563
rect 44545 46523 44603 46529
rect 44818 46520 44824 46572
rect 44876 46560 44882 46572
rect 45189 46563 45247 46569
rect 45189 46560 45201 46563
rect 44876 46532 45201 46560
rect 44876 46520 44882 46532
rect 45189 46529 45201 46532
rect 45235 46529 45247 46563
rect 45830 46560 45836 46572
rect 45791 46532 45836 46560
rect 45189 46523 45247 46529
rect 45830 46520 45836 46532
rect 45888 46520 45894 46572
rect 39482 46492 39488 46504
rect 38436 46464 38700 46492
rect 39443 46464 39488 46492
rect 38436 46452 38442 46464
rect 39482 46452 39488 46464
rect 39540 46452 39546 46504
rect 40678 46492 40684 46504
rect 40639 46464 40684 46492
rect 40678 46452 40684 46464
rect 40736 46452 40742 46504
rect 41506 46452 41512 46504
rect 41564 46492 41570 46504
rect 43901 46495 43959 46501
rect 43901 46492 43913 46495
rect 41564 46464 43913 46492
rect 41564 46452 41570 46464
rect 43901 46461 43913 46464
rect 43947 46461 43959 46495
rect 43901 46455 43959 46461
rect 37366 46424 37372 46436
rect 36464 46396 37372 46424
rect 37366 46384 37372 46396
rect 37424 46384 37430 46436
rect 41325 46427 41383 46433
rect 41325 46424 41337 46427
rect 38580 46396 41337 46424
rect 33100 46328 34468 46356
rect 33100 46316 33106 46328
rect 35618 46316 35624 46368
rect 35676 46356 35682 46368
rect 38580 46356 38608 46396
rect 41325 46393 41337 46396
rect 41371 46393 41383 46427
rect 42613 46427 42671 46433
rect 42613 46424 42625 46427
rect 41325 46387 41383 46393
rect 41432 46396 42625 46424
rect 35676 46328 38608 46356
rect 35676 46316 35682 46328
rect 38930 46316 38936 46368
rect 38988 46356 38994 46368
rect 41432 46356 41460 46396
rect 42613 46393 42625 46396
rect 42659 46393 42671 46427
rect 42613 46387 42671 46393
rect 38988 46328 41460 46356
rect 38988 46316 38994 46328
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 11698 46112 11704 46164
rect 11756 46152 11762 46164
rect 16945 46155 17003 46161
rect 16945 46152 16957 46155
rect 11756 46124 16957 46152
rect 11756 46112 11762 46124
rect 16945 46121 16957 46124
rect 16991 46121 17003 46155
rect 16945 46115 17003 46121
rect 17586 46112 17592 46164
rect 17644 46152 17650 46164
rect 18690 46152 18696 46164
rect 17644 46124 18184 46152
rect 18651 46124 18696 46152
rect 17644 46112 17650 46124
rect 16114 46044 16120 46096
rect 16172 46084 16178 46096
rect 18156 46084 18184 46124
rect 18690 46112 18696 46124
rect 18748 46112 18754 46164
rect 19521 46155 19579 46161
rect 19521 46121 19533 46155
rect 19567 46152 19579 46155
rect 19567 46124 24808 46152
rect 19567 46121 19579 46124
rect 19521 46115 19579 46121
rect 24780 46096 24808 46124
rect 24854 46112 24860 46164
rect 24912 46152 24918 46164
rect 27062 46152 27068 46164
rect 24912 46124 27068 46152
rect 24912 46112 24918 46124
rect 27062 46112 27068 46124
rect 27120 46112 27126 46164
rect 27249 46155 27307 46161
rect 27249 46121 27261 46155
rect 27295 46152 27307 46155
rect 27706 46152 27712 46164
rect 27295 46124 27712 46152
rect 27295 46121 27307 46124
rect 27249 46115 27307 46121
rect 27706 46112 27712 46124
rect 27764 46112 27770 46164
rect 29638 46112 29644 46164
rect 29696 46152 29702 46164
rect 30193 46155 30251 46161
rect 30193 46152 30205 46155
rect 29696 46124 30205 46152
rect 29696 46112 29702 46124
rect 30193 46121 30205 46124
rect 30239 46121 30251 46155
rect 30193 46115 30251 46121
rect 31294 46112 31300 46164
rect 31352 46152 31358 46164
rect 31352 46124 32352 46152
rect 31352 46112 31358 46124
rect 16172 46056 18092 46084
rect 18156 46056 20668 46084
rect 16172 46044 16178 46056
rect 18064 46025 18092 46056
rect 18049 46019 18107 46025
rect 18049 45985 18061 46019
rect 18095 45985 18107 46019
rect 19334 46016 19340 46028
rect 18049 45979 18107 45985
rect 18800 45988 19340 46016
rect 16301 45951 16359 45957
rect 16301 45917 16313 45951
rect 16347 45948 16359 45951
rect 17402 45948 17408 45960
rect 16347 45920 17408 45948
rect 16347 45917 16359 45920
rect 16301 45911 16359 45917
rect 17402 45908 17408 45920
rect 17460 45908 17466 45960
rect 17497 45951 17555 45957
rect 17497 45917 17509 45951
rect 17543 45917 17555 45951
rect 17497 45911 17555 45917
rect 17957 45951 18015 45957
rect 17957 45917 17969 45951
rect 18003 45948 18015 45951
rect 18800 45948 18828 45988
rect 19334 45976 19340 45988
rect 19392 45976 19398 46028
rect 20640 46016 20668 46056
rect 21174 46044 21180 46096
rect 21232 46084 21238 46096
rect 24762 46084 24768 46096
rect 21232 46056 22416 46084
rect 24675 46056 24768 46084
rect 21232 46044 21238 46056
rect 22388 46025 22416 46056
rect 24762 46044 24768 46056
rect 24820 46084 24826 46096
rect 29362 46084 29368 46096
rect 24820 46056 25452 46084
rect 24820 46044 24826 46056
rect 21453 46019 21511 46025
rect 21453 46016 21465 46019
rect 20640 45988 21465 46016
rect 21453 45985 21465 45988
rect 21499 45985 21511 46019
rect 21453 45979 21511 45985
rect 22373 46019 22431 46025
rect 22373 45985 22385 46019
rect 22419 45985 22431 46019
rect 22373 45979 22431 45985
rect 23385 46019 23443 46025
rect 23385 45985 23397 46019
rect 23431 46016 23443 46019
rect 24302 46016 24308 46028
rect 23431 45988 24308 46016
rect 23431 45985 23443 45988
rect 23385 45979 23443 45985
rect 24302 45976 24308 45988
rect 24360 45976 24366 46028
rect 25424 46016 25452 46056
rect 27816 46056 29368 46084
rect 26142 46016 26148 46028
rect 25424 45988 26148 46016
rect 18003 45920 18828 45948
rect 18877 45951 18935 45957
rect 18003 45917 18015 45920
rect 17957 45911 18015 45917
rect 18877 45917 18889 45951
rect 18923 45948 18935 45951
rect 19794 45948 19800 45960
rect 18923 45920 19800 45948
rect 18923 45917 18935 45920
rect 18877 45911 18935 45917
rect 12802 45840 12808 45892
rect 12860 45880 12866 45892
rect 17512 45880 17540 45911
rect 19794 45908 19800 45920
rect 19852 45908 19858 45960
rect 19886 45908 19892 45960
rect 19944 45948 19950 45960
rect 19981 45951 20039 45957
rect 19981 45948 19993 45951
rect 19944 45920 19993 45948
rect 19944 45908 19950 45920
rect 19981 45917 19993 45920
rect 20027 45917 20039 45951
rect 19981 45911 20039 45917
rect 20093 45951 20151 45957
rect 20093 45917 20105 45951
rect 20139 45948 20151 45951
rect 21726 45948 21732 45960
rect 20139 45920 21220 45948
rect 21687 45920 21732 45948
rect 20139 45917 20151 45920
rect 20093 45911 20151 45917
rect 20180 45880 20208 45920
rect 12860 45852 17448 45880
rect 17512 45852 20208 45880
rect 20533 45883 20591 45889
rect 12860 45840 12866 45852
rect 17420 45812 17448 45852
rect 20533 45849 20545 45883
rect 20579 45880 20591 45883
rect 21082 45880 21088 45892
rect 20579 45852 21088 45880
rect 20579 45849 20591 45852
rect 20533 45843 20591 45849
rect 21082 45840 21088 45852
rect 21140 45840 21146 45892
rect 19426 45812 19432 45824
rect 17420 45784 19432 45812
rect 19426 45772 19432 45784
rect 19484 45772 19490 45824
rect 19886 45772 19892 45824
rect 19944 45812 19950 45824
rect 20622 45812 20628 45824
rect 19944 45784 20628 45812
rect 19944 45772 19950 45784
rect 20622 45772 20628 45784
rect 20680 45772 20686 45824
rect 21192 45812 21220 45920
rect 21726 45908 21732 45920
rect 21784 45908 21790 45960
rect 21818 45908 21824 45960
rect 21876 45957 21882 45960
rect 21876 45948 21883 45957
rect 22465 45951 22523 45957
rect 21876 45920 21921 45948
rect 21876 45911 21883 45920
rect 22465 45917 22477 45951
rect 22511 45948 22523 45951
rect 22738 45948 22744 45960
rect 22511 45920 22744 45948
rect 22511 45917 22523 45920
rect 22465 45911 22523 45917
rect 21876 45908 21882 45911
rect 22738 45908 22744 45920
rect 22796 45908 22802 45960
rect 23198 45908 23204 45960
rect 23256 45948 23262 45960
rect 25424 45957 25452 45988
rect 26142 45976 26148 45988
rect 26200 45976 26206 46028
rect 23293 45951 23351 45957
rect 23293 45948 23305 45951
rect 23256 45920 23305 45948
rect 23256 45908 23262 45920
rect 23293 45917 23305 45920
rect 23339 45917 23351 45951
rect 23293 45911 23351 45917
rect 23569 45951 23627 45957
rect 23569 45917 23581 45951
rect 23615 45917 23627 45951
rect 23569 45911 23627 45917
rect 25041 45951 25099 45957
rect 25041 45917 25053 45951
rect 25087 45917 25099 45951
rect 25041 45911 25099 45917
rect 25409 45951 25467 45957
rect 25409 45917 25421 45951
rect 25455 45917 25467 45951
rect 25409 45911 25467 45917
rect 25501 45951 25559 45957
rect 25501 45917 25513 45951
rect 25547 45948 25559 45951
rect 26050 45948 26056 45960
rect 25547 45920 26056 45948
rect 25547 45917 25559 45920
rect 25501 45911 25559 45917
rect 23106 45840 23112 45892
rect 23164 45880 23170 45892
rect 23584 45880 23612 45911
rect 24578 45880 24584 45892
rect 23164 45852 23612 45880
rect 24539 45852 24584 45880
rect 23164 45840 23170 45852
rect 24578 45840 24584 45852
rect 24636 45840 24642 45892
rect 25056 45880 25084 45911
rect 26050 45908 26056 45920
rect 26108 45908 26114 45960
rect 26234 45948 26240 45960
rect 26195 45920 26240 45948
rect 26234 45908 26240 45920
rect 26292 45908 26298 45960
rect 26326 45908 26332 45960
rect 26384 45948 26390 45960
rect 26789 45951 26847 45957
rect 26384 45920 26429 45948
rect 26384 45908 26390 45920
rect 26789 45917 26801 45951
rect 26835 45917 26847 45951
rect 26789 45911 26847 45917
rect 26344 45880 26372 45908
rect 25056 45852 26372 45880
rect 26418 45840 26424 45892
rect 26476 45880 26482 45892
rect 26804 45880 26832 45911
rect 26970 45908 26976 45960
rect 27028 45948 27034 45960
rect 27816 45948 27844 46056
rect 29362 46044 29368 46056
rect 29420 46044 29426 46096
rect 30926 46044 30932 46096
rect 30984 46084 30990 46096
rect 31665 46087 31723 46093
rect 31665 46084 31677 46087
rect 30984 46056 31677 46084
rect 30984 46044 30990 46056
rect 31665 46053 31677 46056
rect 31711 46053 31723 46087
rect 31665 46047 31723 46053
rect 32324 46084 32352 46124
rect 33226 46112 33232 46164
rect 33284 46152 33290 46164
rect 34330 46152 34336 46164
rect 33284 46124 34336 46152
rect 33284 46112 33290 46124
rect 34330 46112 34336 46124
rect 34388 46152 34394 46164
rect 35710 46152 35716 46164
rect 34388 46124 35716 46152
rect 34388 46112 34394 46124
rect 35710 46112 35716 46124
rect 35768 46112 35774 46164
rect 36354 46152 36360 46164
rect 36315 46124 36360 46152
rect 36354 46112 36360 46124
rect 36412 46112 36418 46164
rect 39298 46112 39304 46164
rect 39356 46152 39362 46164
rect 42337 46155 42395 46161
rect 42337 46152 42349 46155
rect 39356 46124 42349 46152
rect 39356 46112 39362 46124
rect 42337 46121 42349 46124
rect 42383 46121 42395 46155
rect 42337 46115 42395 46121
rect 42610 46112 42616 46164
rect 42668 46152 42674 46164
rect 43625 46155 43683 46161
rect 43625 46152 43637 46155
rect 42668 46124 43637 46152
rect 42668 46112 42674 46124
rect 43625 46121 43637 46124
rect 43671 46121 43683 46155
rect 44266 46152 44272 46164
rect 44227 46124 44272 46152
rect 43625 46115 43683 46121
rect 44266 46112 44272 46124
rect 44324 46112 44330 46164
rect 32324 46056 40632 46084
rect 27890 45976 27896 46028
rect 27948 46016 27954 46028
rect 27948 45988 30972 46016
rect 32324 46002 32352 46056
rect 33045 46019 33103 46025
rect 27948 45976 27954 45988
rect 28902 45948 28908 45960
rect 27028 45920 27844 45948
rect 28863 45920 28908 45948
rect 27028 45908 27034 45920
rect 28902 45908 28908 45920
rect 28960 45908 28966 45960
rect 29181 45951 29239 45957
rect 29181 45917 29193 45951
rect 29227 45917 29239 45951
rect 29181 45911 29239 45917
rect 26476 45852 26832 45880
rect 26476 45840 26482 45852
rect 27614 45840 27620 45892
rect 27672 45880 27678 45892
rect 28445 45883 28503 45889
rect 28445 45880 28457 45883
rect 27672 45852 28457 45880
rect 27672 45840 27678 45852
rect 28445 45849 28457 45852
rect 28491 45849 28503 45883
rect 28994 45880 29000 45892
rect 28955 45852 29000 45880
rect 28445 45843 28503 45849
rect 28994 45840 29000 45852
rect 29052 45840 29058 45892
rect 29196 45880 29224 45911
rect 29362 45908 29368 45960
rect 29420 45948 29426 45960
rect 29733 45951 29791 45957
rect 29733 45948 29745 45951
rect 29420 45920 29745 45948
rect 29420 45908 29426 45920
rect 29733 45917 29745 45920
rect 29779 45948 29791 45951
rect 29822 45948 29828 45960
rect 29779 45920 29828 45948
rect 29779 45917 29791 45920
rect 29733 45911 29791 45917
rect 29822 45908 29828 45920
rect 29880 45908 29886 45960
rect 30101 45951 30159 45957
rect 30101 45917 30113 45951
rect 30147 45948 30159 45951
rect 30282 45948 30288 45960
rect 30147 45920 30288 45948
rect 30147 45917 30159 45920
rect 30101 45911 30159 45917
rect 30282 45908 30288 45920
rect 30340 45908 30346 45960
rect 30944 45957 30972 45988
rect 33045 45985 33057 46019
rect 33091 46016 33103 46019
rect 33134 46016 33140 46028
rect 33091 45988 33140 46016
rect 33091 45985 33103 45988
rect 33045 45979 33103 45985
rect 33134 45976 33140 45988
rect 33192 45976 33198 46028
rect 33502 45976 33508 46028
rect 33560 46016 33566 46028
rect 36832 46025 36860 46056
rect 40604 46028 40632 46056
rect 41138 46044 41144 46096
rect 41196 46084 41202 46096
rect 42981 46087 43039 46093
rect 42981 46084 42993 46087
rect 41196 46056 42993 46084
rect 41196 46044 41202 46056
rect 42981 46053 42993 46056
rect 43027 46053 43039 46087
rect 42981 46047 43039 46053
rect 35529 46019 35587 46025
rect 35529 46016 35541 46019
rect 33560 45988 35541 46016
rect 33560 45976 33566 45988
rect 35529 45985 35541 45988
rect 35575 45985 35587 46019
rect 35529 45979 35587 45985
rect 36817 46019 36875 46025
rect 36817 45985 36829 46019
rect 36863 45985 36875 46019
rect 37550 46016 37556 46028
rect 36817 45979 36875 45985
rect 37292 45988 37556 46016
rect 30929 45951 30987 45957
rect 30929 45917 30941 45951
rect 30975 45917 30987 45951
rect 32030 45948 32036 45960
rect 31991 45920 32036 45948
rect 30929 45911 30987 45917
rect 32030 45908 32036 45920
rect 32088 45908 32094 45960
rect 32677 45951 32735 45957
rect 32677 45917 32689 45951
rect 32723 45948 32735 45951
rect 33410 45948 33416 45960
rect 32723 45920 33416 45948
rect 32723 45917 32735 45920
rect 32677 45911 32735 45917
rect 33410 45908 33416 45920
rect 33468 45948 33474 45960
rect 33686 45948 33692 45960
rect 33468 45920 33692 45948
rect 33468 45908 33474 45920
rect 33686 45908 33692 45920
rect 33744 45908 33750 45960
rect 33870 45948 33876 45960
rect 33831 45920 33876 45948
rect 33870 45908 33876 45920
rect 33928 45908 33934 45960
rect 34885 45951 34943 45957
rect 34885 45948 34897 45951
rect 34164 45920 34897 45948
rect 30190 45880 30196 45892
rect 29196 45852 30196 45880
rect 30190 45840 30196 45852
rect 30248 45840 30254 45892
rect 31938 45840 31944 45892
rect 31996 45880 32002 45892
rect 33505 45883 33563 45889
rect 33505 45880 33517 45883
rect 31996 45852 33517 45880
rect 31996 45840 32002 45852
rect 33505 45849 33517 45852
rect 33551 45849 33563 45883
rect 34054 45880 34060 45892
rect 34015 45852 34060 45880
rect 33505 45843 33563 45849
rect 34054 45840 34060 45852
rect 34112 45840 34118 45892
rect 25406 45812 25412 45824
rect 21192 45784 25412 45812
rect 25406 45772 25412 45784
rect 25464 45772 25470 45824
rect 27798 45772 27804 45824
rect 27856 45812 27862 45824
rect 27893 45815 27951 45821
rect 27893 45812 27905 45815
rect 27856 45784 27905 45812
rect 27856 45772 27862 45784
rect 27893 45781 27905 45784
rect 27939 45781 27951 45815
rect 27893 45775 27951 45781
rect 31478 45772 31484 45824
rect 31536 45812 31542 45824
rect 34164 45812 34192 45920
rect 34885 45917 34897 45920
rect 34931 45917 34943 45951
rect 36906 45948 36912 45960
rect 36867 45920 36912 45948
rect 34885 45911 34943 45917
rect 36906 45908 36912 45920
rect 36964 45908 36970 45960
rect 37292 45957 37320 45988
rect 37550 45976 37556 45988
rect 37608 46016 37614 46028
rect 38470 46016 38476 46028
rect 37608 45988 38476 46016
rect 37608 45976 37614 45988
rect 38470 45976 38476 45988
rect 38528 45976 38534 46028
rect 39209 46019 39267 46025
rect 39209 45985 39221 46019
rect 39255 46016 39267 46019
rect 39482 46016 39488 46028
rect 39255 45988 39488 46016
rect 39255 45985 39267 45988
rect 39209 45979 39267 45985
rect 39482 45976 39488 45988
rect 39540 45976 39546 46028
rect 40586 46016 40592 46028
rect 40547 45988 40592 46016
rect 40586 45976 40592 45988
rect 40644 45976 40650 46028
rect 42242 45976 42248 46028
rect 42300 46016 42306 46028
rect 44284 46016 44312 46112
rect 42300 45988 44312 46016
rect 42300 45976 42306 45988
rect 37277 45951 37335 45957
rect 37277 45917 37289 45951
rect 37323 45917 37335 45951
rect 37277 45911 37335 45917
rect 37461 45951 37519 45957
rect 37461 45917 37473 45951
rect 37507 45948 37519 45951
rect 37642 45948 37648 45960
rect 37507 45920 37648 45948
rect 37507 45917 37519 45920
rect 37461 45911 37519 45917
rect 37642 45908 37648 45920
rect 37700 45908 37706 45960
rect 38289 45951 38347 45957
rect 38289 45917 38301 45951
rect 38335 45948 38347 45951
rect 38562 45948 38568 45960
rect 38335 45920 38568 45948
rect 38335 45917 38347 45920
rect 38289 45911 38347 45917
rect 38562 45908 38568 45920
rect 38620 45908 38626 45960
rect 39114 45948 39120 45960
rect 39075 45920 39120 45948
rect 39114 45908 39120 45920
rect 39172 45908 39178 45960
rect 39574 45908 39580 45960
rect 39632 45948 39638 45960
rect 40681 45951 40739 45957
rect 40681 45948 40693 45951
rect 39632 45920 40693 45948
rect 39632 45908 39638 45920
rect 40681 45917 40693 45920
rect 40727 45917 40739 45951
rect 40681 45911 40739 45917
rect 34422 45840 34428 45892
rect 34480 45880 34486 45892
rect 38102 45880 38108 45892
rect 34480 45852 38108 45880
rect 34480 45840 34486 45852
rect 38102 45840 38108 45852
rect 38160 45840 38166 45892
rect 38194 45840 38200 45892
rect 38252 45880 38258 45892
rect 38381 45883 38439 45889
rect 38381 45880 38393 45883
rect 38252 45852 38393 45880
rect 38252 45840 38258 45852
rect 38381 45849 38393 45852
rect 38427 45849 38439 45883
rect 38580 45880 38608 45908
rect 40126 45880 40132 45892
rect 38580 45852 40132 45880
rect 38381 45843 38439 45849
rect 40126 45840 40132 45852
rect 40184 45840 40190 45892
rect 40696 45880 40724 45911
rect 40770 45908 40776 45960
rect 40828 45948 40834 45960
rect 41141 45951 41199 45957
rect 41141 45948 41153 45951
rect 40828 45920 41153 45948
rect 40828 45908 40834 45920
rect 41141 45917 41153 45920
rect 41187 45917 41199 45951
rect 41141 45911 41199 45917
rect 41230 45908 41236 45960
rect 41288 45948 41294 45960
rect 41288 45920 41333 45948
rect 41288 45908 41294 45920
rect 42242 45880 42248 45892
rect 40696 45852 42248 45880
rect 42242 45840 42248 45852
rect 42300 45840 42306 45892
rect 31536 45784 34192 45812
rect 31536 45772 31542 45784
rect 41414 45772 41420 45824
rect 41472 45812 41478 45824
rect 41693 45815 41751 45821
rect 41693 45812 41705 45815
rect 41472 45784 41705 45812
rect 41472 45772 41478 45784
rect 41693 45781 41705 45784
rect 41739 45781 41751 45815
rect 41693 45775 41751 45781
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 17126 45568 17132 45620
rect 17184 45608 17190 45620
rect 17184 45580 19012 45608
rect 17184 45568 17190 45580
rect 18984 45484 19012 45580
rect 19334 45568 19340 45620
rect 19392 45608 19398 45620
rect 20530 45608 20536 45620
rect 19392 45580 20536 45608
rect 19392 45568 19398 45580
rect 20530 45568 20536 45580
rect 20588 45568 20594 45620
rect 20622 45568 20628 45620
rect 20680 45608 20686 45620
rect 23661 45611 23719 45617
rect 20680 45580 22508 45608
rect 20680 45568 20686 45580
rect 17865 45475 17923 45481
rect 17865 45441 17877 45475
rect 17911 45472 17923 45475
rect 17954 45472 17960 45484
rect 17911 45444 17960 45472
rect 17911 45441 17923 45444
rect 17865 45435 17923 45441
rect 17954 45432 17960 45444
rect 18012 45432 18018 45484
rect 18782 45472 18788 45484
rect 18743 45444 18788 45472
rect 18782 45432 18788 45444
rect 18840 45432 18846 45484
rect 18966 45432 18972 45484
rect 19024 45472 19030 45484
rect 19337 45475 19395 45481
rect 19024 45444 19117 45472
rect 19024 45432 19030 45444
rect 19337 45441 19349 45475
rect 19383 45472 19395 45475
rect 20533 45475 20591 45481
rect 20533 45472 20545 45475
rect 19383 45444 20545 45472
rect 19383 45441 19395 45444
rect 19337 45435 19395 45441
rect 20533 45441 20545 45444
rect 20579 45441 20591 45475
rect 20898 45472 20904 45484
rect 20859 45444 20904 45472
rect 20533 45435 20591 45441
rect 20898 45432 20904 45444
rect 20956 45432 20962 45484
rect 20990 45432 20996 45484
rect 21048 45472 21054 45484
rect 22480 45481 22508 45580
rect 23661 45577 23673 45611
rect 23707 45608 23719 45611
rect 23842 45608 23848 45620
rect 23707 45580 23848 45608
rect 23707 45577 23719 45580
rect 23661 45571 23719 45577
rect 23842 45568 23848 45580
rect 23900 45568 23906 45620
rect 24302 45568 24308 45620
rect 24360 45608 24366 45620
rect 27522 45608 27528 45620
rect 24360 45580 27528 45608
rect 24360 45568 24366 45580
rect 27522 45568 27528 45580
rect 27580 45568 27586 45620
rect 29270 45568 29276 45620
rect 29328 45608 29334 45620
rect 29328 45580 31524 45608
rect 29328 45568 29334 45580
rect 23474 45540 23480 45552
rect 22848 45512 23480 45540
rect 22848 45481 22876 45512
rect 23474 45500 23480 45512
rect 23532 45540 23538 45552
rect 24578 45540 24584 45552
rect 23532 45512 24584 45540
rect 23532 45500 23538 45512
rect 24578 45500 24584 45512
rect 24636 45500 24642 45552
rect 24857 45543 24915 45549
rect 24857 45509 24869 45543
rect 24903 45540 24915 45543
rect 25130 45540 25136 45552
rect 24903 45512 25136 45540
rect 24903 45509 24915 45512
rect 24857 45503 24915 45509
rect 25130 45500 25136 45512
rect 25188 45500 25194 45552
rect 25314 45500 25320 45552
rect 25372 45540 25378 45552
rect 25372 45512 28212 45540
rect 25372 45500 25378 45512
rect 21085 45475 21143 45481
rect 21085 45472 21097 45475
rect 21048 45444 21097 45472
rect 21048 45432 21054 45444
rect 21085 45441 21097 45444
rect 21131 45472 21143 45475
rect 22465 45475 22523 45481
rect 21131 45444 22094 45472
rect 21131 45441 21143 45444
rect 21085 45435 21143 45441
rect 4614 45364 4620 45416
rect 4672 45404 4678 45416
rect 18325 45407 18383 45413
rect 18325 45404 18337 45407
rect 4672 45376 18337 45404
rect 4672 45364 4678 45376
rect 18325 45373 18337 45376
rect 18371 45373 18383 45407
rect 18325 45367 18383 45373
rect 19245 45407 19303 45413
rect 19245 45373 19257 45407
rect 19291 45404 19303 45407
rect 20162 45404 20168 45416
rect 19291 45376 20168 45404
rect 19291 45373 19303 45376
rect 19245 45367 19303 45373
rect 20162 45364 20168 45376
rect 20220 45364 20226 45416
rect 17221 45339 17279 45345
rect 17221 45305 17233 45339
rect 17267 45336 17279 45339
rect 20622 45336 20628 45348
rect 17267 45308 20628 45336
rect 17267 45305 17279 45308
rect 17221 45299 17279 45305
rect 20622 45296 20628 45308
rect 20680 45296 20686 45348
rect 22066 45336 22094 45444
rect 22465 45441 22477 45475
rect 22511 45441 22523 45475
rect 22465 45435 22523 45441
rect 22833 45475 22891 45481
rect 22833 45441 22845 45475
rect 22879 45441 22891 45475
rect 23198 45472 23204 45484
rect 23159 45444 23204 45472
rect 22833 45435 22891 45441
rect 23198 45432 23204 45444
rect 23256 45432 23262 45484
rect 25406 45432 25412 45484
rect 25464 45472 25470 45484
rect 25501 45475 25559 45481
rect 25501 45472 25513 45475
rect 25464 45444 25513 45472
rect 25464 45432 25470 45444
rect 25501 45441 25513 45444
rect 25547 45441 25559 45475
rect 25501 45435 25559 45441
rect 25869 45475 25927 45481
rect 25869 45441 25881 45475
rect 25915 45441 25927 45475
rect 26050 45472 26056 45484
rect 26011 45444 26056 45472
rect 25869 45435 25927 45441
rect 22925 45407 22983 45413
rect 22925 45373 22937 45407
rect 22971 45404 22983 45407
rect 23014 45404 23020 45416
rect 22971 45376 23020 45404
rect 22971 45373 22983 45376
rect 22925 45367 22983 45373
rect 23014 45364 23020 45376
rect 23072 45364 23078 45416
rect 23106 45364 23112 45416
rect 23164 45404 23170 45416
rect 25593 45407 25651 45413
rect 23164 45376 23209 45404
rect 23164 45364 23170 45376
rect 25593 45373 25605 45407
rect 25639 45373 25651 45407
rect 25884 45404 25912 45435
rect 26050 45432 26056 45444
rect 26108 45432 26114 45484
rect 26142 45432 26148 45484
rect 26200 45472 26206 45484
rect 28184 45481 28212 45512
rect 29932 45512 31064 45540
rect 29932 45484 29960 45512
rect 31036 45484 31064 45512
rect 26513 45475 26571 45481
rect 26513 45472 26525 45475
rect 26200 45444 26525 45472
rect 26200 45432 26206 45444
rect 26513 45441 26525 45444
rect 26559 45441 26571 45475
rect 26513 45435 26571 45441
rect 28169 45475 28227 45481
rect 28169 45441 28181 45475
rect 28215 45441 28227 45475
rect 28169 45435 28227 45441
rect 28537 45475 28595 45481
rect 28537 45441 28549 45475
rect 28583 45441 28595 45475
rect 28537 45435 28595 45441
rect 28629 45475 28687 45481
rect 28629 45441 28641 45475
rect 28675 45472 28687 45475
rect 28902 45472 28908 45484
rect 28675 45444 28908 45472
rect 28675 45441 28687 45444
rect 28629 45435 28687 45441
rect 26418 45404 26424 45416
rect 25884 45376 26424 45404
rect 25593 45367 25651 45373
rect 25498 45336 25504 45348
rect 22066 45308 25504 45336
rect 25498 45296 25504 45308
rect 25556 45296 25562 45348
rect 25608 45336 25636 45367
rect 26418 45364 26424 45376
rect 26476 45404 26482 45416
rect 28442 45404 28448 45416
rect 26476 45376 28448 45404
rect 26476 45364 26482 45376
rect 28442 45364 28448 45376
rect 28500 45364 28506 45416
rect 28552 45404 28580 45435
rect 28902 45432 28908 45444
rect 28960 45472 28966 45484
rect 29365 45475 29423 45481
rect 29365 45472 29377 45475
rect 28960 45444 29377 45472
rect 28960 45432 28966 45444
rect 29365 45441 29377 45444
rect 29411 45441 29423 45475
rect 29914 45472 29920 45484
rect 29365 45435 29423 45441
rect 29656 45444 29920 45472
rect 28994 45404 29000 45416
rect 28552 45376 29000 45404
rect 28994 45364 29000 45376
rect 29052 45364 29058 45416
rect 29273 45407 29331 45413
rect 29273 45373 29285 45407
rect 29319 45404 29331 45407
rect 29656 45404 29684 45444
rect 29914 45432 29920 45444
rect 29972 45432 29978 45484
rect 30006 45432 30012 45484
rect 30064 45472 30070 45484
rect 30101 45475 30159 45481
rect 30101 45472 30113 45475
rect 30064 45444 30113 45472
rect 30064 45432 30070 45444
rect 30101 45441 30113 45444
rect 30147 45441 30159 45475
rect 31018 45472 31024 45484
rect 30931 45444 31024 45472
rect 30101 45435 30159 45441
rect 31018 45432 31024 45444
rect 31076 45432 31082 45484
rect 31496 45481 31524 45580
rect 36262 45568 36268 45620
rect 36320 45608 36326 45620
rect 40586 45608 40592 45620
rect 36320 45580 40592 45608
rect 36320 45568 36326 45580
rect 40586 45568 40592 45580
rect 40644 45608 40650 45620
rect 41230 45608 41236 45620
rect 40644 45580 41236 45608
rect 40644 45568 40650 45580
rect 41230 45568 41236 45580
rect 41288 45568 41294 45620
rect 43898 45608 43904 45620
rect 43811 45580 43904 45608
rect 43898 45568 43904 45580
rect 43956 45608 43962 45620
rect 45186 45608 45192 45620
rect 43956 45580 45192 45608
rect 43956 45568 43962 45580
rect 45186 45568 45192 45580
rect 45244 45568 45250 45620
rect 34701 45543 34759 45549
rect 34701 45509 34713 45543
rect 34747 45540 34759 45543
rect 34790 45540 34796 45552
rect 34747 45512 34796 45540
rect 34747 45509 34759 45512
rect 34701 45503 34759 45509
rect 34790 45500 34796 45512
rect 34848 45500 34854 45552
rect 35618 45540 35624 45552
rect 34900 45512 35624 45540
rect 31481 45475 31539 45481
rect 31481 45441 31493 45475
rect 31527 45441 31539 45475
rect 31481 45435 31539 45441
rect 33042 45432 33048 45484
rect 33100 45472 33106 45484
rect 33321 45475 33379 45481
rect 33321 45472 33333 45475
rect 33100 45444 33333 45472
rect 33100 45432 33106 45444
rect 33321 45441 33333 45444
rect 33367 45472 33379 45475
rect 33410 45472 33416 45484
rect 33367 45444 33416 45472
rect 33367 45441 33379 45444
rect 33321 45435 33379 45441
rect 33410 45432 33416 45444
rect 33468 45432 33474 45484
rect 33689 45475 33747 45481
rect 33689 45441 33701 45475
rect 33735 45472 33747 45475
rect 34900 45472 34928 45512
rect 35618 45500 35624 45512
rect 35676 45540 35682 45552
rect 35713 45543 35771 45549
rect 35713 45540 35725 45543
rect 35676 45512 35725 45540
rect 35676 45500 35682 45512
rect 35713 45509 35725 45512
rect 35759 45509 35771 45543
rect 35713 45503 35771 45509
rect 36630 45500 36636 45552
rect 36688 45540 36694 45552
rect 40681 45543 40739 45549
rect 40681 45540 40693 45543
rect 36688 45512 40693 45540
rect 36688 45500 36694 45512
rect 40681 45509 40693 45512
rect 40727 45540 40739 45543
rect 41782 45540 41788 45552
rect 40727 45512 41788 45540
rect 40727 45509 40739 45512
rect 40681 45503 40739 45509
rect 41782 45500 41788 45512
rect 41840 45500 41846 45552
rect 33735 45444 34928 45472
rect 35069 45475 35127 45481
rect 33735 45441 33747 45444
rect 33689 45435 33747 45441
rect 35069 45441 35081 45475
rect 35115 45441 35127 45475
rect 35069 45435 35127 45441
rect 35253 45475 35311 45481
rect 35253 45441 35265 45475
rect 35299 45472 35311 45475
rect 36449 45475 36507 45481
rect 35299 45444 35756 45472
rect 35299 45441 35311 45444
rect 35253 45435 35311 45441
rect 29319 45376 29684 45404
rect 29319 45373 29331 45376
rect 29273 45367 29331 45373
rect 29730 45364 29736 45416
rect 29788 45404 29794 45416
rect 30193 45407 30251 45413
rect 30193 45404 30205 45407
rect 29788 45376 30205 45404
rect 29788 45364 29794 45376
rect 30193 45373 30205 45376
rect 30239 45373 30251 45407
rect 34054 45404 34060 45416
rect 34015 45376 34060 45404
rect 30193 45367 30251 45373
rect 34054 45364 34060 45376
rect 34112 45364 34118 45416
rect 35084 45404 35112 45435
rect 35728 45416 35756 45444
rect 36449 45441 36461 45475
rect 36495 45441 36507 45475
rect 36722 45472 36728 45484
rect 36683 45444 36728 45472
rect 36449 45435 36507 45441
rect 35526 45404 35532 45416
rect 35084 45376 35532 45404
rect 35526 45364 35532 45376
rect 35584 45364 35590 45416
rect 35710 45364 35716 45416
rect 35768 45364 35774 45416
rect 36262 45404 36268 45416
rect 36223 45376 36268 45404
rect 36262 45364 36268 45376
rect 36320 45364 36326 45416
rect 26326 45336 26332 45348
rect 25608 45308 26332 45336
rect 26326 45296 26332 45308
rect 26384 45296 26390 45348
rect 26602 45336 26608 45348
rect 26436 45308 26608 45336
rect 20073 45271 20131 45277
rect 20073 45237 20085 45271
rect 20119 45268 20131 45271
rect 24210 45268 24216 45280
rect 20119 45240 24216 45268
rect 20119 45237 20131 45240
rect 20073 45231 20131 45237
rect 24210 45228 24216 45240
rect 24268 45228 24274 45280
rect 24397 45271 24455 45277
rect 24397 45237 24409 45271
rect 24443 45268 24455 45271
rect 25222 45268 25228 45280
rect 24443 45240 25228 45268
rect 24443 45237 24455 45240
rect 24397 45231 24455 45237
rect 25222 45228 25228 45240
rect 25280 45268 25286 45280
rect 26436 45268 26464 45308
rect 26602 45296 26608 45308
rect 26660 45296 26666 45348
rect 27982 45336 27988 45348
rect 27943 45308 27988 45336
rect 27982 45296 27988 45308
rect 28040 45296 28046 45348
rect 28460 45336 28488 45364
rect 30374 45336 30380 45348
rect 28460 45308 30380 45336
rect 30374 45296 30380 45308
rect 30432 45336 30438 45348
rect 30837 45339 30895 45345
rect 30837 45336 30849 45339
rect 30432 45308 30849 45336
rect 30432 45296 30438 45308
rect 30837 45305 30849 45308
rect 30883 45305 30895 45339
rect 36464 45336 36492 45435
rect 36722 45432 36728 45444
rect 36780 45432 36786 45484
rect 38102 45472 38108 45484
rect 38063 45444 38108 45472
rect 38102 45432 38108 45444
rect 38160 45432 38166 45484
rect 38473 45475 38531 45481
rect 38473 45441 38485 45475
rect 38519 45472 38531 45475
rect 38654 45472 38660 45484
rect 38519 45444 38660 45472
rect 38519 45441 38531 45444
rect 38473 45435 38531 45441
rect 38654 45432 38660 45444
rect 38712 45432 38718 45484
rect 39114 45472 39120 45484
rect 39027 45444 39120 45472
rect 39114 45432 39120 45444
rect 39172 45432 39178 45484
rect 40310 45472 40316 45484
rect 40271 45444 40316 45472
rect 40310 45432 40316 45444
rect 40368 45432 40374 45484
rect 40770 45472 40776 45484
rect 40683 45444 40776 45472
rect 40770 45432 40776 45444
rect 40828 45432 40834 45484
rect 41506 45472 41512 45484
rect 41467 45444 41512 45472
rect 41506 45432 41512 45444
rect 41564 45432 41570 45484
rect 42610 45472 42616 45484
rect 42571 45444 42616 45472
rect 42610 45432 42616 45444
rect 42668 45432 42674 45484
rect 36909 45407 36967 45413
rect 36909 45373 36921 45407
rect 36955 45404 36967 45407
rect 37182 45404 37188 45416
rect 36955 45376 37188 45404
rect 36955 45373 36967 45376
rect 36909 45367 36967 45373
rect 37182 45364 37188 45376
rect 37240 45404 37246 45416
rect 37642 45404 37648 45416
rect 37240 45376 37648 45404
rect 37240 45364 37246 45376
rect 37642 45364 37648 45376
rect 37700 45364 37706 45416
rect 38194 45364 38200 45416
rect 38252 45404 38258 45416
rect 38562 45404 38568 45416
rect 38252 45376 38568 45404
rect 38252 45364 38258 45376
rect 38562 45364 38568 45376
rect 38620 45364 38626 45416
rect 39132 45404 39160 45432
rect 40402 45404 40408 45416
rect 39132 45376 40408 45404
rect 37366 45336 37372 45348
rect 36464 45308 37372 45336
rect 30837 45299 30895 45305
rect 37366 45296 37372 45308
rect 37424 45336 37430 45348
rect 37550 45336 37556 45348
rect 37424 45308 37556 45336
rect 37424 45296 37430 45308
rect 37550 45296 37556 45308
rect 37608 45296 37614 45348
rect 37921 45339 37979 45345
rect 37921 45305 37933 45339
rect 37967 45336 37979 45339
rect 38286 45336 38292 45348
rect 37967 45308 38292 45336
rect 37967 45305 37979 45308
rect 37921 45299 37979 45305
rect 38286 45296 38292 45308
rect 38344 45296 38350 45348
rect 27246 45268 27252 45280
rect 25280 45240 26464 45268
rect 27207 45240 27252 45268
rect 25280 45228 25286 45240
rect 27246 45228 27252 45240
rect 27304 45228 27310 45280
rect 27798 45228 27804 45280
rect 27856 45268 27862 45280
rect 29546 45268 29552 45280
rect 27856 45240 29552 45268
rect 27856 45228 27862 45240
rect 29546 45228 29552 45240
rect 29604 45228 29610 45280
rect 37642 45228 37648 45280
rect 37700 45268 37706 45280
rect 39132 45268 39160 45376
rect 40402 45364 40408 45376
rect 40460 45364 40466 45416
rect 40586 45404 40592 45416
rect 40547 45376 40592 45404
rect 40586 45364 40592 45376
rect 40644 45364 40650 45416
rect 39850 45336 39856 45348
rect 39811 45308 39856 45336
rect 39850 45296 39856 45308
rect 39908 45296 39914 45348
rect 39298 45268 39304 45280
rect 37700 45240 39160 45268
rect 39259 45240 39304 45268
rect 37700 45228 37706 45240
rect 39298 45228 39304 45240
rect 39356 45268 39362 45280
rect 40788 45268 40816 45432
rect 43254 45364 43260 45416
rect 43312 45404 43318 45416
rect 43809 45407 43867 45413
rect 43809 45404 43821 45407
rect 43312 45376 43821 45404
rect 43312 45364 43318 45376
rect 43809 45373 43821 45376
rect 43855 45404 43867 45407
rect 43916 45404 43944 45568
rect 43855 45376 43944 45404
rect 43855 45373 43867 45376
rect 43809 45367 43867 45373
rect 39356 45240 40816 45268
rect 39356 45228 39362 45240
rect 42702 45228 42708 45280
rect 42760 45268 42766 45280
rect 43257 45271 43315 45277
rect 43257 45268 43269 45271
rect 42760 45240 43269 45268
rect 42760 45228 42766 45240
rect 43257 45237 43269 45240
rect 43303 45237 43315 45271
rect 43257 45231 43315 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 18322 45064 18328 45076
rect 18283 45036 18328 45064
rect 18322 45024 18328 45036
rect 18380 45024 18386 45076
rect 24029 45067 24087 45073
rect 24029 45033 24041 45067
rect 24075 45064 24087 45067
rect 24946 45064 24952 45076
rect 24075 45036 24952 45064
rect 24075 45033 24087 45036
rect 24029 45027 24087 45033
rect 24946 45024 24952 45036
rect 25004 45024 25010 45076
rect 25498 45024 25504 45076
rect 25556 45064 25562 45076
rect 34146 45064 34152 45076
rect 25556 45036 31156 45064
rect 34107 45036 34152 45064
rect 25556 45024 25562 45036
rect 23106 44956 23112 45008
rect 23164 44996 23170 45008
rect 24857 44999 24915 45005
rect 24857 44996 24869 44999
rect 23164 44968 24869 44996
rect 23164 44956 23170 44968
rect 24857 44965 24869 44968
rect 24903 44996 24915 44999
rect 25590 44996 25596 45008
rect 24903 44968 25596 44996
rect 24903 44965 24915 44968
rect 24857 44959 24915 44965
rect 25590 44956 25596 44968
rect 25648 44956 25654 45008
rect 26050 44956 26056 45008
rect 26108 44996 26114 45008
rect 28721 44999 28779 45005
rect 28721 44996 28733 44999
rect 26108 44968 28733 44996
rect 26108 44956 26114 44968
rect 28721 44965 28733 44968
rect 28767 44965 28779 44999
rect 28721 44959 28779 44965
rect 29730 44956 29736 45008
rect 29788 44996 29794 45008
rect 31128 45005 31156 45036
rect 34146 45024 34152 45036
rect 34204 45024 34210 45076
rect 39942 45024 39948 45076
rect 40000 45064 40006 45076
rect 40037 45067 40095 45073
rect 40037 45064 40049 45067
rect 40000 45036 40049 45064
rect 40000 45024 40006 45036
rect 40037 45033 40049 45036
rect 40083 45033 40095 45067
rect 42242 45064 42248 45076
rect 42203 45036 42248 45064
rect 40037 45027 40095 45033
rect 42242 45024 42248 45036
rect 42300 45024 42306 45076
rect 30009 44999 30067 45005
rect 30009 44996 30021 44999
rect 29788 44968 30021 44996
rect 29788 44956 29794 44968
rect 30009 44965 30021 44968
rect 30055 44965 30067 44999
rect 30009 44959 30067 44965
rect 31113 44999 31171 45005
rect 31113 44965 31125 44999
rect 31159 44965 31171 44999
rect 34974 44996 34980 45008
rect 31113 44959 31171 44965
rect 31220 44968 34980 44996
rect 20625 44931 20683 44937
rect 20625 44897 20637 44931
rect 20671 44928 20683 44931
rect 20898 44928 20904 44940
rect 20671 44900 20904 44928
rect 20671 44897 20683 44900
rect 20625 44891 20683 44897
rect 20898 44888 20904 44900
rect 20956 44928 20962 44940
rect 23385 44931 23443 44937
rect 20956 44900 23152 44928
rect 20956 44888 20962 44900
rect 18138 44860 18144 44872
rect 18099 44832 18144 44860
rect 18138 44820 18144 44832
rect 18196 44820 18202 44872
rect 19978 44860 19984 44872
rect 19939 44832 19984 44860
rect 19978 44820 19984 44832
rect 20036 44820 20042 44872
rect 20533 44863 20591 44869
rect 20533 44829 20545 44863
rect 20579 44860 20591 44863
rect 20990 44860 20996 44872
rect 20579 44832 20996 44860
rect 20579 44829 20591 44832
rect 20533 44823 20591 44829
rect 20990 44820 20996 44832
rect 21048 44820 21054 44872
rect 22002 44860 22008 44872
rect 21963 44832 22008 44860
rect 22002 44820 22008 44832
rect 22060 44820 22066 44872
rect 22925 44863 22983 44869
rect 22925 44829 22937 44863
rect 22971 44860 22983 44863
rect 23014 44860 23020 44872
rect 22971 44832 23020 44860
rect 22971 44829 22983 44832
rect 22925 44823 22983 44829
rect 23014 44820 23020 44832
rect 23072 44820 23078 44872
rect 22186 44792 22192 44804
rect 22147 44764 22192 44792
rect 22186 44752 22192 44764
rect 22244 44752 22250 44804
rect 23124 44792 23152 44900
rect 23385 44897 23397 44931
rect 23431 44928 23443 44931
rect 24118 44928 24124 44940
rect 23431 44900 24124 44928
rect 23431 44897 23443 44900
rect 23385 44891 23443 44897
rect 24118 44888 24124 44900
rect 24176 44888 24182 44940
rect 25406 44928 25412 44940
rect 25367 44900 25412 44928
rect 25406 44888 25412 44900
rect 25464 44888 25470 44940
rect 28077 44931 28135 44937
rect 26252 44900 27844 44928
rect 26252 44872 26280 44900
rect 23201 44863 23259 44869
rect 23201 44829 23213 44863
rect 23247 44860 23259 44863
rect 23474 44860 23480 44872
rect 23247 44832 23480 44860
rect 23247 44829 23259 44832
rect 23201 44823 23259 44829
rect 23474 44820 23480 44832
rect 23532 44820 23538 44872
rect 24210 44820 24216 44872
rect 24268 44860 24274 44872
rect 24673 44863 24731 44869
rect 24673 44860 24685 44863
rect 24268 44832 24685 44860
rect 24268 44820 24274 44832
rect 24673 44829 24685 44832
rect 24719 44829 24731 44863
rect 24673 44823 24731 44829
rect 25314 44820 25320 44872
rect 25372 44860 25378 44872
rect 25958 44860 25964 44872
rect 25372 44832 25964 44860
rect 25372 44820 25378 44832
rect 25958 44820 25964 44832
rect 26016 44820 26022 44872
rect 26234 44860 26240 44872
rect 26195 44832 26240 44860
rect 26234 44820 26240 44832
rect 26292 44820 26298 44872
rect 26418 44860 26424 44872
rect 26379 44832 26424 44860
rect 26418 44820 26424 44832
rect 26476 44820 26482 44872
rect 27614 44860 27620 44872
rect 27575 44832 27620 44860
rect 27614 44820 27620 44832
rect 27672 44820 27678 44872
rect 27154 44792 27160 44804
rect 23124 44764 24992 44792
rect 27115 44764 27160 44792
rect 18782 44684 18788 44736
rect 18840 44724 18846 44736
rect 19797 44727 19855 44733
rect 19797 44724 19809 44727
rect 18840 44696 19809 44724
rect 18840 44684 18846 44696
rect 19797 44693 19809 44696
rect 19843 44693 19855 44727
rect 21910 44724 21916 44736
rect 21871 44696 21916 44724
rect 19797 44687 19855 44693
rect 21910 44684 21916 44696
rect 21968 44684 21974 44736
rect 22370 44684 22376 44736
rect 22428 44724 22434 44736
rect 24302 44724 24308 44736
rect 22428 44696 24308 44724
rect 22428 44684 22434 44696
rect 24302 44684 24308 44696
rect 24360 44684 24366 44736
rect 24964 44724 24992 44764
rect 27154 44752 27160 44764
rect 27212 44752 27218 44804
rect 27816 44792 27844 44900
rect 28077 44897 28089 44931
rect 28123 44928 28135 44931
rect 29638 44928 29644 44940
rect 28123 44900 29644 44928
rect 28123 44897 28135 44900
rect 28077 44891 28135 44897
rect 29638 44888 29644 44900
rect 29696 44888 29702 44940
rect 30282 44888 30288 44940
rect 30340 44928 30346 44940
rect 31220 44928 31248 44968
rect 34974 44956 34980 44968
rect 35032 44956 35038 45008
rect 35161 44999 35219 45005
rect 35161 44965 35173 44999
rect 35207 44996 35219 44999
rect 35342 44996 35348 45008
rect 35207 44968 35348 44996
rect 35207 44965 35219 44968
rect 35161 44959 35219 44965
rect 35342 44956 35348 44968
rect 35400 44956 35406 45008
rect 33410 44928 33416 44940
rect 30340 44900 31248 44928
rect 31726 44900 33416 44928
rect 30340 44888 30346 44900
rect 27982 44860 27988 44872
rect 27943 44832 27988 44860
rect 27982 44820 27988 44832
rect 28040 44820 28046 44872
rect 28905 44863 28963 44869
rect 28905 44829 28917 44863
rect 28951 44829 28963 44863
rect 28905 44823 28963 44829
rect 28920 44792 28948 44823
rect 29546 44820 29552 44872
rect 29604 44860 29610 44872
rect 29733 44863 29791 44869
rect 29733 44860 29745 44863
rect 29604 44832 29745 44860
rect 29604 44820 29610 44832
rect 29733 44829 29745 44832
rect 29779 44829 29791 44863
rect 29733 44823 29791 44829
rect 30377 44863 30435 44869
rect 30377 44829 30389 44863
rect 30423 44860 30435 44863
rect 31726 44860 31754 44900
rect 33410 44888 33416 44900
rect 33468 44888 33474 44940
rect 34054 44928 34060 44940
rect 33612 44900 34060 44928
rect 31938 44860 31944 44872
rect 30423 44832 31754 44860
rect 31899 44832 31944 44860
rect 30423 44829 30435 44832
rect 30377 44823 30435 44829
rect 30392 44792 30420 44823
rect 31938 44820 31944 44832
rect 31996 44820 32002 44872
rect 32030 44820 32036 44872
rect 32088 44860 32094 44872
rect 32306 44860 32312 44872
rect 32088 44832 32133 44860
rect 32267 44832 32312 44860
rect 32088 44820 32094 44832
rect 32306 44820 32312 44832
rect 32364 44820 32370 44872
rect 33612 44869 33640 44900
rect 34054 44888 34060 44900
rect 34112 44888 34118 44940
rect 36262 44888 36268 44940
rect 36320 44928 36326 44940
rect 37001 44931 37059 44937
rect 37001 44928 37013 44931
rect 36320 44900 37013 44928
rect 36320 44888 36326 44900
rect 37001 44897 37013 44900
rect 37047 44928 37059 44931
rect 39482 44928 39488 44940
rect 37047 44900 39488 44928
rect 37047 44897 37059 44900
rect 37001 44891 37059 44897
rect 33597 44863 33655 44869
rect 33597 44829 33609 44863
rect 33643 44829 33655 44863
rect 33597 44823 33655 44829
rect 33689 44863 33747 44869
rect 33689 44829 33701 44863
rect 33735 44860 33747 44863
rect 33962 44860 33968 44872
rect 33735 44832 33968 44860
rect 33735 44829 33747 44832
rect 33689 44823 33747 44829
rect 33962 44820 33968 44832
rect 34020 44820 34026 44872
rect 34885 44863 34943 44869
rect 34885 44829 34897 44863
rect 34931 44829 34943 44863
rect 35526 44860 35532 44872
rect 35487 44832 35532 44860
rect 34885 44823 34943 44829
rect 27816 44764 30420 44792
rect 31573 44795 31631 44801
rect 31573 44761 31585 44795
rect 31619 44792 31631 44795
rect 33134 44792 33140 44804
rect 31619 44764 31754 44792
rect 33095 44764 33140 44792
rect 31619 44761 31631 44764
rect 31573 44755 31631 44761
rect 28166 44724 28172 44736
rect 24964 44696 28172 44724
rect 28166 44684 28172 44696
rect 28224 44684 28230 44736
rect 31726 44724 31754 44764
rect 33134 44752 33140 44764
rect 33192 44752 33198 44804
rect 34606 44724 34612 44736
rect 31726 44696 34612 44724
rect 34606 44684 34612 44696
rect 34664 44724 34670 44736
rect 34900 44724 34928 44823
rect 35526 44820 35532 44832
rect 35584 44820 35590 44872
rect 35710 44860 35716 44872
rect 35671 44832 35716 44860
rect 35710 44820 35716 44832
rect 35768 44820 35774 44872
rect 37277 44863 37335 44869
rect 37277 44829 37289 44863
rect 37323 44860 37335 44863
rect 37366 44860 37372 44872
rect 37323 44832 37372 44860
rect 37323 44829 37335 44832
rect 37277 44823 37335 44829
rect 37366 44820 37372 44832
rect 37424 44820 37430 44872
rect 37461 44863 37519 44869
rect 37461 44829 37473 44863
rect 37507 44860 37519 44863
rect 37550 44860 37556 44872
rect 37507 44832 37556 44860
rect 37507 44829 37519 44832
rect 37461 44823 37519 44829
rect 37550 44820 37556 44832
rect 37608 44820 37614 44872
rect 38197 44863 38255 44869
rect 38197 44829 38209 44863
rect 38243 44829 38255 44863
rect 38654 44860 38660 44872
rect 38615 44832 38660 44860
rect 38197 44823 38255 44829
rect 36446 44792 36452 44804
rect 36407 44764 36452 44792
rect 36446 44752 36452 44764
rect 36504 44752 36510 44804
rect 37384 44792 37412 44820
rect 38212 44792 38240 44823
rect 38654 44820 38660 44832
rect 38712 44820 38718 44872
rect 38948 44869 38976 44900
rect 39482 44888 39488 44900
rect 39540 44888 39546 44940
rect 40310 44888 40316 44940
rect 40368 44928 40374 44940
rect 40681 44931 40739 44937
rect 40681 44928 40693 44931
rect 40368 44900 40693 44928
rect 40368 44888 40374 44900
rect 40681 44897 40693 44900
rect 40727 44897 40739 44931
rect 40681 44891 40739 44897
rect 41233 44931 41291 44937
rect 41233 44897 41245 44931
rect 41279 44928 41291 44931
rect 41414 44928 41420 44940
rect 41279 44900 41420 44928
rect 41279 44897 41291 44900
rect 41233 44891 41291 44897
rect 41414 44888 41420 44900
rect 41472 44888 41478 44940
rect 42702 44928 42708 44940
rect 41524 44900 42708 44928
rect 38933 44863 38991 44869
rect 38933 44829 38945 44863
rect 38979 44829 38991 44863
rect 39298 44860 39304 44872
rect 39259 44832 39304 44860
rect 38933 44823 38991 44829
rect 39298 44820 39304 44832
rect 39356 44820 39362 44872
rect 41322 44820 41328 44872
rect 41380 44860 41386 44872
rect 41524 44869 41552 44900
rect 42702 44888 42708 44900
rect 42760 44888 42766 44940
rect 41509 44863 41567 44869
rect 41509 44860 41521 44863
rect 41380 44832 41521 44860
rect 41380 44820 41386 44832
rect 41509 44829 41521 44832
rect 41555 44829 41567 44863
rect 41509 44823 41567 44829
rect 41693 44863 41751 44869
rect 41693 44829 41705 44863
rect 41739 44829 41751 44863
rect 41693 44823 41751 44829
rect 37384 44764 38240 44792
rect 40770 44752 40776 44804
rect 40828 44792 40834 44804
rect 41708 44792 41736 44823
rect 40828 44764 41736 44792
rect 40828 44752 40834 44764
rect 34664 44696 34928 44724
rect 34664 44684 34670 44696
rect 36170 44684 36176 44736
rect 36228 44724 36234 44736
rect 37182 44724 37188 44736
rect 36228 44696 37188 44724
rect 36228 44684 36234 44696
rect 37182 44684 37188 44696
rect 37240 44724 37246 44736
rect 40218 44724 40224 44736
rect 37240 44696 40224 44724
rect 37240 44684 37246 44696
rect 40218 44684 40224 44696
rect 40276 44684 40282 44736
rect 43254 44724 43260 44736
rect 43215 44696 43260 44724
rect 43254 44684 43260 44696
rect 43312 44684 43318 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 18966 44480 18972 44532
rect 19024 44520 19030 44532
rect 19613 44523 19671 44529
rect 19613 44520 19625 44523
rect 19024 44492 19625 44520
rect 19024 44480 19030 44492
rect 19613 44489 19625 44492
rect 19659 44489 19671 44523
rect 19613 44483 19671 44489
rect 20530 44480 20536 44532
rect 20588 44520 20594 44532
rect 21269 44523 21327 44529
rect 21269 44520 21281 44523
rect 20588 44492 21281 44520
rect 20588 44480 20594 44492
rect 21269 44489 21281 44492
rect 21315 44489 21327 44523
rect 21269 44483 21327 44489
rect 22002 44480 22008 44532
rect 22060 44520 22066 44532
rect 22370 44520 22376 44532
rect 22060 44492 22376 44520
rect 22060 44480 22066 44492
rect 22370 44480 22376 44492
rect 22428 44480 22434 44532
rect 23106 44520 23112 44532
rect 22756 44492 23112 44520
rect 18046 44412 18052 44464
rect 18104 44452 18110 44464
rect 18325 44455 18383 44461
rect 18325 44452 18337 44455
rect 18104 44424 18337 44452
rect 18104 44412 18110 44424
rect 18325 44421 18337 44424
rect 18371 44452 18383 44455
rect 18371 44424 21220 44452
rect 18371 44421 18383 44424
rect 18325 44415 18383 44421
rect 19058 44384 19064 44396
rect 19019 44356 19064 44384
rect 19058 44344 19064 44356
rect 19116 44344 19122 44396
rect 19797 44387 19855 44393
rect 19797 44353 19809 44387
rect 19843 44384 19855 44387
rect 19978 44384 19984 44396
rect 19843 44356 19984 44384
rect 19843 44353 19855 44356
rect 19797 44347 19855 44353
rect 19978 44344 19984 44356
rect 20036 44344 20042 44396
rect 20349 44387 20407 44393
rect 20349 44353 20361 44387
rect 20395 44353 20407 44387
rect 20530 44384 20536 44396
rect 20491 44356 20536 44384
rect 20349 44347 20407 44353
rect 20364 44316 20392 44347
rect 20530 44344 20536 44356
rect 20588 44344 20594 44396
rect 21082 44384 21088 44396
rect 21043 44356 21088 44384
rect 21082 44344 21088 44356
rect 21140 44344 21146 44396
rect 21192 44384 21220 44424
rect 21910 44412 21916 44464
rect 21968 44452 21974 44464
rect 22646 44452 22652 44464
rect 21968 44424 22652 44452
rect 21968 44412 21974 44424
rect 22646 44412 22652 44424
rect 22704 44412 22710 44464
rect 22465 44387 22523 44393
rect 21192 44356 22416 44384
rect 20714 44316 20720 44328
rect 20364 44288 20720 44316
rect 20714 44276 20720 44288
rect 20772 44316 20778 44328
rect 22005 44319 22063 44325
rect 22005 44316 22017 44319
rect 20772 44288 22017 44316
rect 20772 44276 20778 44288
rect 22005 44285 22017 44288
rect 22051 44285 22063 44319
rect 22005 44279 22063 44285
rect 22388 44248 22416 44356
rect 22465 44353 22477 44387
rect 22511 44384 22523 44387
rect 22756 44384 22784 44492
rect 23106 44480 23112 44492
rect 23164 44480 23170 44532
rect 24210 44480 24216 44532
rect 24268 44520 24274 44532
rect 26326 44520 26332 44532
rect 24268 44492 26188 44520
rect 26287 44492 26332 44520
rect 24268 44480 24274 44492
rect 22830 44412 22836 44464
rect 22888 44452 22894 44464
rect 22888 44424 22933 44452
rect 22888 44412 22894 44424
rect 23014 44412 23020 44464
rect 23072 44452 23078 44464
rect 23753 44455 23811 44461
rect 23753 44452 23765 44455
rect 23072 44424 23765 44452
rect 23072 44412 23078 44424
rect 23753 44421 23765 44424
rect 23799 44421 23811 44455
rect 26160 44452 26188 44492
rect 26326 44480 26332 44492
rect 26384 44480 26390 44532
rect 27798 44520 27804 44532
rect 27356 44492 27804 44520
rect 27356 44452 27384 44492
rect 27798 44480 27804 44492
rect 27856 44480 27862 44532
rect 39850 44520 39856 44532
rect 28092 44492 39856 44520
rect 27982 44452 27988 44464
rect 23753 44415 23811 44421
rect 24596 44424 25452 44452
rect 22922 44384 22928 44396
rect 22511 44356 22784 44384
rect 22883 44356 22928 44384
rect 22511 44353 22523 44356
rect 22465 44347 22523 44353
rect 22922 44344 22928 44356
rect 22980 44344 22986 44396
rect 24302 44384 24308 44396
rect 24263 44356 24308 44384
rect 24302 44344 24308 44356
rect 24360 44344 24366 44396
rect 24596 44393 24624 44424
rect 24581 44387 24639 44393
rect 24581 44353 24593 44387
rect 24627 44353 24639 44387
rect 24762 44384 24768 44396
rect 24723 44356 24768 44384
rect 24581 44347 24639 44353
rect 24762 44344 24768 44356
rect 24820 44344 24826 44396
rect 25222 44384 25228 44396
rect 25183 44356 25228 44384
rect 25222 44344 25228 44356
rect 25280 44344 25286 44396
rect 25424 44393 25452 44424
rect 26160 44424 27384 44452
rect 27448 44424 27988 44452
rect 25409 44387 25467 44393
rect 25409 44353 25421 44387
rect 25455 44384 25467 44387
rect 26050 44384 26056 44396
rect 25455 44356 26056 44384
rect 25455 44353 25467 44356
rect 25409 44347 25467 44353
rect 26050 44344 26056 44356
rect 26108 44344 26114 44396
rect 26160 44384 26188 44424
rect 27448 44393 27476 44424
rect 27982 44412 27988 44424
rect 28040 44412 28046 44464
rect 26329 44387 26387 44393
rect 26329 44384 26341 44387
rect 26160 44356 26341 44384
rect 26329 44353 26341 44356
rect 26375 44353 26387 44387
rect 26329 44347 26387 44353
rect 27433 44387 27491 44393
rect 27433 44353 27445 44387
rect 27479 44353 27491 44387
rect 27433 44347 27491 44353
rect 27614 44344 27620 44396
rect 27672 44384 27678 44396
rect 27801 44387 27859 44393
rect 27801 44384 27813 44387
rect 27672 44356 27813 44384
rect 27672 44344 27678 44356
rect 27801 44353 27813 44356
rect 27847 44353 27859 44387
rect 27801 44347 27859 44353
rect 23106 44316 23112 44328
rect 23067 44288 23112 44316
rect 23106 44276 23112 44288
rect 23164 44276 23170 44328
rect 25777 44319 25835 44325
rect 25777 44285 25789 44319
rect 25823 44316 25835 44319
rect 27338 44316 27344 44328
rect 25823 44288 27344 44316
rect 25823 44285 25835 44288
rect 25777 44279 25835 44285
rect 27338 44276 27344 44288
rect 27396 44276 27402 44328
rect 28092 44248 28120 44492
rect 39850 44480 39856 44492
rect 39908 44480 39914 44532
rect 41322 44480 41328 44532
rect 41380 44520 41386 44532
rect 41877 44523 41935 44529
rect 41877 44520 41889 44523
rect 41380 44492 41889 44520
rect 41380 44480 41386 44492
rect 41877 44489 41889 44492
rect 41923 44489 41935 44523
rect 41877 44483 41935 44489
rect 42242 44480 42248 44532
rect 42300 44520 42306 44532
rect 42613 44523 42671 44529
rect 42613 44520 42625 44523
rect 42300 44492 42625 44520
rect 42300 44480 42306 44492
rect 42613 44489 42625 44492
rect 42659 44489 42671 44523
rect 42613 44483 42671 44489
rect 28169 44455 28227 44461
rect 28169 44421 28181 44455
rect 28215 44452 28227 44455
rect 29086 44452 29092 44464
rect 28215 44424 29092 44452
rect 28215 44421 28227 44424
rect 28169 44415 28227 44421
rect 29086 44412 29092 44424
rect 29144 44412 29150 44464
rect 33410 44452 33416 44464
rect 31220 44424 31984 44452
rect 33371 44424 33416 44452
rect 28442 44344 28448 44396
rect 28500 44384 28506 44396
rect 28721 44387 28779 44393
rect 28721 44384 28733 44387
rect 28500 44356 28733 44384
rect 28500 44344 28506 44356
rect 28721 44353 28733 44356
rect 28767 44353 28779 44387
rect 28721 44347 28779 44353
rect 29457 44387 29515 44393
rect 29457 44353 29469 44387
rect 29503 44353 29515 44387
rect 29822 44384 29828 44396
rect 29783 44356 29828 44384
rect 29457 44347 29515 44353
rect 28994 44316 29000 44328
rect 28955 44288 29000 44316
rect 28994 44276 29000 44288
rect 29052 44276 29058 44328
rect 29472 44316 29500 44347
rect 29822 44344 29828 44356
rect 29880 44344 29886 44396
rect 31220 44393 31248 44424
rect 31956 44396 31984 44424
rect 33410 44412 33416 44424
rect 33468 44452 33474 44464
rect 34422 44452 34428 44464
rect 33468 44424 34428 44452
rect 33468 44412 33474 44424
rect 34422 44412 34428 44424
rect 34480 44412 34486 44464
rect 34974 44452 34980 44464
rect 34935 44424 34980 44452
rect 34974 44412 34980 44424
rect 35032 44412 35038 44464
rect 38120 44424 39988 44452
rect 31205 44387 31263 44393
rect 31205 44353 31217 44387
rect 31251 44353 31263 44387
rect 31205 44347 31263 44353
rect 31573 44387 31631 44393
rect 31573 44353 31585 44387
rect 31619 44384 31631 44387
rect 31619 44356 31754 44384
rect 31619 44353 31631 44356
rect 31573 44347 31631 44353
rect 29730 44316 29736 44328
rect 29472 44288 29736 44316
rect 29730 44276 29736 44288
rect 29788 44276 29794 44328
rect 30929 44319 30987 44325
rect 30929 44285 30941 44319
rect 30975 44316 30987 44319
rect 30975 44288 31616 44316
rect 30975 44285 30987 44288
rect 30929 44279 30987 44285
rect 31588 44260 31616 44288
rect 22388 44220 28120 44248
rect 28166 44208 28172 44260
rect 28224 44248 28230 44260
rect 31481 44251 31539 44257
rect 31481 44248 31493 44251
rect 28224 44220 31493 44248
rect 28224 44208 28230 44220
rect 31481 44217 31493 44220
rect 31527 44217 31539 44251
rect 31481 44211 31539 44217
rect 31570 44208 31576 44260
rect 31628 44208 31634 44260
rect 31726 44180 31754 44356
rect 31938 44344 31944 44396
rect 31996 44384 32002 44396
rect 32401 44387 32459 44393
rect 32401 44384 32413 44387
rect 31996 44356 32413 44384
rect 31996 44344 32002 44356
rect 32401 44353 32413 44356
rect 32447 44353 32459 44387
rect 34330 44384 34336 44396
rect 34291 44356 34336 44384
rect 32401 44347 32459 44353
rect 34330 44344 34336 44356
rect 34388 44344 34394 44396
rect 34517 44387 34575 44393
rect 34517 44353 34529 44387
rect 34563 44384 34575 44387
rect 34606 44384 34612 44396
rect 34563 44356 34612 44384
rect 34563 44353 34575 44356
rect 34517 44347 34575 44353
rect 34606 44344 34612 44356
rect 34664 44344 34670 44396
rect 35618 44384 35624 44396
rect 35579 44356 35624 44384
rect 35618 44344 35624 44356
rect 35676 44344 35682 44396
rect 36170 44384 36176 44396
rect 36131 44356 36176 44384
rect 36170 44344 36176 44356
rect 36228 44344 36234 44396
rect 38120 44393 38148 44424
rect 37461 44387 37519 44393
rect 37461 44384 37473 44387
rect 36280 44356 37473 44384
rect 31846 44276 31852 44328
rect 31904 44316 31910 44328
rect 32769 44319 32827 44325
rect 32769 44316 32781 44319
rect 31904 44288 32781 44316
rect 31904 44276 31910 44288
rect 32769 44285 32781 44288
rect 32815 44285 32827 44319
rect 32769 44279 32827 44285
rect 32861 44319 32919 44325
rect 32861 44285 32873 44319
rect 32907 44316 32919 44319
rect 33134 44316 33140 44328
rect 32907 44288 33140 44316
rect 32907 44285 32919 44288
rect 32861 44279 32919 44285
rect 33134 44276 33140 44288
rect 33192 44316 33198 44328
rect 33686 44316 33692 44328
rect 33192 44288 33692 44316
rect 33192 44276 33198 44288
rect 33686 44276 33692 44288
rect 33744 44276 33750 44328
rect 34790 44276 34796 44328
rect 34848 44316 34854 44328
rect 35710 44316 35716 44328
rect 34848 44288 35716 44316
rect 34848 44276 34854 44288
rect 35710 44276 35716 44288
rect 35768 44316 35774 44328
rect 36280 44316 36308 44356
rect 37461 44353 37473 44356
rect 37507 44353 37519 44387
rect 37461 44347 37519 44353
rect 37921 44387 37979 44393
rect 37921 44353 37933 44387
rect 37967 44353 37979 44387
rect 37921 44347 37979 44353
rect 38105 44387 38163 44393
rect 38105 44353 38117 44387
rect 38151 44353 38163 44387
rect 38286 44384 38292 44396
rect 38247 44356 38292 44384
rect 38105 44347 38163 44353
rect 35768 44288 36308 44316
rect 35768 44276 35774 44288
rect 36354 44276 36360 44328
rect 36412 44316 36418 44328
rect 36412 44288 36457 44316
rect 36412 44276 36418 44288
rect 35621 44251 35679 44257
rect 35621 44248 35633 44251
rect 32416 44220 35633 44248
rect 32030 44180 32036 44192
rect 31726 44152 32036 44180
rect 32030 44140 32036 44152
rect 32088 44180 32094 44192
rect 32416 44180 32444 44220
rect 35621 44217 35633 44220
rect 35667 44217 35679 44251
rect 37936 44248 37964 44347
rect 38286 44344 38292 44356
rect 38344 44384 38350 44396
rect 38933 44387 38991 44393
rect 38933 44384 38945 44387
rect 38344 44356 38945 44384
rect 38344 44344 38350 44356
rect 38933 44353 38945 44356
rect 38979 44353 38991 44387
rect 38933 44347 38991 44353
rect 39301 44387 39359 44393
rect 39301 44353 39313 44387
rect 39347 44353 39359 44387
rect 39301 44347 39359 44353
rect 38470 44276 38476 44328
rect 38528 44316 38534 44328
rect 39316 44316 39344 44347
rect 39960 44328 39988 44424
rect 40402 44412 40408 44464
rect 40460 44452 40466 44464
rect 41417 44455 41475 44461
rect 41417 44452 41429 44455
rect 40460 44424 41429 44452
rect 40460 44412 40466 44424
rect 41417 44421 41429 44424
rect 41463 44421 41475 44455
rect 41417 44415 41475 44421
rect 40497 44387 40555 44393
rect 40497 44353 40509 44387
rect 40543 44384 40555 44387
rect 40586 44384 40592 44396
rect 40543 44356 40592 44384
rect 40543 44353 40555 44356
rect 40497 44347 40555 44353
rect 40586 44344 40592 44356
rect 40644 44344 40650 44396
rect 40770 44344 40776 44396
rect 40828 44384 40834 44396
rect 40865 44387 40923 44393
rect 40865 44384 40877 44387
rect 40828 44356 40877 44384
rect 40828 44344 40834 44356
rect 40865 44353 40877 44356
rect 40911 44353 40923 44387
rect 40865 44347 40923 44353
rect 38528 44288 39344 44316
rect 38528 44276 38534 44288
rect 39942 44276 39948 44328
rect 40000 44316 40006 44328
rect 40129 44319 40187 44325
rect 40129 44316 40141 44319
rect 40000 44288 40141 44316
rect 40000 44276 40006 44288
rect 40129 44285 40141 44288
rect 40175 44285 40187 44319
rect 40129 44279 40187 44285
rect 38488 44248 38516 44276
rect 41874 44248 41880 44260
rect 37936 44220 38516 44248
rect 38856 44220 41880 44248
rect 35621 44211 35679 44217
rect 32088 44152 32444 44180
rect 32088 44140 32094 44152
rect 34146 44140 34152 44192
rect 34204 44180 34210 44192
rect 34241 44183 34299 44189
rect 34241 44180 34253 44183
rect 34204 44152 34253 44180
rect 34204 44140 34210 44152
rect 34241 44149 34253 44152
rect 34287 44149 34299 44183
rect 34241 44143 34299 44149
rect 34422 44140 34428 44192
rect 34480 44180 34486 44192
rect 38856 44180 38884 44220
rect 41874 44208 41880 44220
rect 41932 44208 41938 44260
rect 39390 44180 39396 44192
rect 34480 44152 38884 44180
rect 39351 44152 39396 44180
rect 34480 44140 34486 44152
rect 39390 44140 39396 44152
rect 39448 44140 39454 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 21726 43936 21732 43988
rect 21784 43976 21790 43988
rect 24029 43979 24087 43985
rect 21784 43948 22140 43976
rect 21784 43936 21790 43948
rect 20530 43868 20536 43920
rect 20588 43908 20594 43920
rect 22005 43911 22063 43917
rect 22005 43908 22017 43911
rect 20588 43880 22017 43908
rect 20588 43868 20594 43880
rect 22005 43877 22017 43880
rect 22051 43877 22063 43911
rect 22112 43908 22140 43948
rect 24029 43945 24041 43979
rect 24075 43976 24087 43979
rect 24394 43976 24400 43988
rect 24075 43948 24400 43976
rect 24075 43945 24087 43948
rect 24029 43939 24087 43945
rect 24394 43936 24400 43948
rect 24452 43936 24458 43988
rect 28258 43936 28264 43988
rect 28316 43976 28322 43988
rect 28905 43979 28963 43985
rect 28905 43976 28917 43979
rect 28316 43948 28917 43976
rect 28316 43936 28322 43948
rect 28905 43945 28917 43948
rect 28951 43945 28963 43979
rect 30098 43976 30104 43988
rect 30059 43948 30104 43976
rect 28905 43939 28963 43945
rect 30098 43936 30104 43948
rect 30156 43936 30162 43988
rect 31110 43976 31116 43988
rect 31071 43948 31116 43976
rect 31110 43936 31116 43948
rect 31168 43936 31174 43988
rect 31754 43936 31760 43988
rect 31812 43976 31818 43988
rect 32306 43976 32312 43988
rect 31812 43948 32312 43976
rect 31812 43936 31818 43948
rect 32306 43936 32312 43948
rect 32364 43976 32370 43988
rect 33229 43979 33287 43985
rect 33229 43976 33241 43979
rect 32364 43948 33241 43976
rect 32364 43936 32370 43948
rect 33229 43945 33241 43948
rect 33275 43945 33287 43979
rect 37274 43976 37280 43988
rect 37235 43948 37280 43976
rect 33229 43939 33287 43945
rect 37274 43936 37280 43948
rect 37332 43936 37338 43988
rect 38381 43979 38439 43985
rect 38381 43945 38393 43979
rect 38427 43976 38439 43979
rect 38470 43976 38476 43988
rect 38427 43948 38476 43976
rect 38427 43945 38439 43948
rect 38381 43939 38439 43945
rect 38470 43936 38476 43948
rect 38528 43936 38534 43988
rect 40586 43976 40592 43988
rect 40547 43948 40592 43976
rect 40586 43936 40592 43948
rect 40644 43936 40650 43988
rect 41785 43979 41843 43985
rect 41785 43945 41797 43979
rect 41831 43976 41843 43979
rect 43254 43976 43260 43988
rect 41831 43948 43260 43976
rect 41831 43945 41843 43948
rect 41785 43939 41843 43945
rect 43254 43936 43260 43948
rect 43312 43936 43318 43988
rect 22112 43880 27016 43908
rect 22005 43871 22063 43877
rect 20162 43840 20168 43852
rect 20123 43812 20168 43840
rect 20162 43800 20168 43812
rect 20220 43800 20226 43852
rect 21910 43840 21916 43852
rect 21744 43812 21916 43840
rect 20530 43772 20536 43784
rect 20491 43744 20536 43772
rect 20530 43732 20536 43744
rect 20588 43732 20594 43784
rect 20714 43772 20720 43784
rect 20675 43744 20720 43772
rect 20714 43732 20720 43744
rect 20772 43732 20778 43784
rect 21744 43781 21772 43812
rect 21910 43800 21916 43812
rect 21968 43840 21974 43852
rect 26988 43849 27016 43880
rect 27246 43868 27252 43920
rect 27304 43908 27310 43920
rect 30558 43908 30564 43920
rect 27304 43880 30564 43908
rect 27304 43868 27310 43880
rect 30558 43868 30564 43880
rect 30616 43868 30622 43920
rect 26973 43843 27031 43849
rect 21968 43812 22876 43840
rect 21968 43800 21974 43812
rect 21453 43775 21511 43781
rect 21453 43741 21465 43775
rect 21499 43741 21511 43775
rect 21453 43735 21511 43741
rect 21729 43775 21787 43781
rect 21729 43741 21741 43775
rect 21775 43741 21787 43775
rect 21729 43735 21787 43741
rect 22281 43775 22339 43781
rect 22281 43741 22293 43775
rect 22327 43772 22339 43775
rect 22738 43772 22744 43784
rect 22327 43744 22744 43772
rect 22327 43741 22339 43744
rect 22281 43735 22339 43741
rect 21468 43704 21496 43735
rect 22738 43732 22744 43744
rect 22796 43732 22802 43784
rect 22848 43781 22876 43812
rect 26973 43809 26985 43843
rect 27019 43809 27031 43843
rect 33686 43840 33692 43852
rect 33647 43812 33692 43840
rect 26973 43803 27031 43809
rect 33686 43800 33692 43812
rect 33744 43800 33750 43852
rect 38102 43800 38108 43852
rect 38160 43840 38166 43852
rect 38841 43843 38899 43849
rect 38841 43840 38853 43843
rect 38160 43812 38853 43840
rect 38160 43800 38166 43812
rect 38841 43809 38853 43812
rect 38887 43840 38899 43843
rect 39301 43843 39359 43849
rect 39301 43840 39313 43843
rect 38887 43812 39313 43840
rect 38887 43809 38899 43812
rect 38841 43803 38899 43809
rect 39301 43809 39313 43812
rect 39347 43840 39359 43843
rect 40037 43843 40095 43849
rect 40037 43840 40049 43843
rect 39347 43812 40049 43840
rect 39347 43809 39359 43812
rect 39301 43803 39359 43809
rect 40037 43809 40049 43812
rect 40083 43809 40095 43843
rect 40037 43803 40095 43809
rect 22833 43775 22891 43781
rect 22833 43741 22845 43775
rect 22879 43741 22891 43775
rect 22833 43735 22891 43741
rect 24762 43732 24768 43784
rect 24820 43772 24826 43784
rect 25501 43775 25559 43781
rect 25501 43772 25513 43775
rect 24820 43744 25513 43772
rect 24820 43732 24826 43744
rect 25501 43741 25513 43744
rect 25547 43741 25559 43775
rect 25501 43735 25559 43741
rect 26421 43775 26479 43781
rect 26421 43741 26433 43775
rect 26467 43772 26479 43775
rect 26467 43744 27292 43772
rect 26467 43741 26479 43744
rect 26421 43735 26479 43741
rect 23106 43704 23112 43716
rect 21468 43676 23112 43704
rect 23106 43664 23112 43676
rect 23164 43664 23170 43716
rect 23290 43704 23296 43716
rect 23251 43676 23296 43704
rect 23290 43664 23296 43676
rect 23348 43664 23354 43716
rect 23382 43664 23388 43716
rect 23440 43704 23446 43716
rect 24581 43707 24639 43713
rect 24581 43704 24593 43707
rect 23440 43676 24593 43704
rect 23440 43664 23446 43676
rect 24581 43673 24593 43676
rect 24627 43673 24639 43707
rect 27264 43704 27292 43744
rect 27338 43732 27344 43784
rect 27396 43772 27402 43784
rect 27433 43775 27491 43781
rect 27433 43772 27445 43775
rect 27396 43744 27445 43772
rect 27396 43732 27402 43744
rect 27433 43741 27445 43744
rect 27479 43741 27491 43775
rect 27614 43772 27620 43784
rect 27575 43744 27620 43772
rect 27433 43735 27491 43741
rect 27614 43732 27620 43744
rect 27672 43732 27678 43784
rect 27798 43772 27804 43784
rect 27759 43744 27804 43772
rect 27798 43732 27804 43744
rect 27856 43732 27862 43784
rect 28074 43772 28080 43784
rect 28035 43744 28080 43772
rect 28074 43732 28080 43744
rect 28132 43732 28138 43784
rect 28166 43732 28172 43784
rect 28224 43772 28230 43784
rect 28353 43775 28411 43781
rect 28353 43772 28365 43775
rect 28224 43744 28365 43772
rect 28224 43732 28230 43744
rect 28353 43741 28365 43744
rect 28399 43741 28411 43775
rect 28353 43735 28411 43741
rect 31573 43775 31631 43781
rect 31573 43741 31585 43775
rect 31619 43772 31631 43775
rect 31846 43772 31852 43784
rect 31619 43744 31852 43772
rect 31619 43741 31631 43744
rect 31573 43735 31631 43741
rect 31846 43732 31852 43744
rect 31904 43732 31910 43784
rect 32217 43775 32275 43781
rect 32217 43741 32229 43775
rect 32263 43772 32275 43775
rect 32766 43772 32772 43784
rect 32263 43744 32772 43772
rect 32263 43741 32275 43744
rect 32217 43735 32275 43741
rect 32766 43732 32772 43744
rect 32824 43732 32830 43784
rect 33778 43772 33784 43784
rect 33739 43744 33784 43772
rect 33778 43732 33784 43744
rect 33836 43732 33842 43784
rect 34146 43772 34152 43784
rect 34107 43744 34152 43772
rect 34146 43732 34152 43744
rect 34204 43732 34210 43784
rect 34333 43775 34391 43781
rect 34333 43741 34345 43775
rect 34379 43772 34391 43775
rect 34514 43772 34520 43784
rect 34379 43744 34520 43772
rect 34379 43741 34391 43744
rect 34333 43735 34391 43741
rect 34514 43732 34520 43744
rect 34572 43772 34578 43784
rect 34790 43772 34796 43784
rect 34572 43744 34796 43772
rect 34572 43732 34578 43744
rect 34790 43732 34796 43744
rect 34848 43732 34854 43784
rect 35437 43775 35495 43781
rect 35437 43772 35449 43775
rect 35176 43744 35449 43772
rect 27982 43704 27988 43716
rect 27264 43676 27988 43704
rect 24581 43667 24639 43673
rect 27982 43664 27988 43676
rect 28040 43664 28046 43716
rect 34422 43664 34428 43716
rect 34480 43704 34486 43716
rect 35176 43704 35204 43744
rect 35437 43741 35449 43744
rect 35483 43741 35495 43775
rect 35437 43735 35495 43741
rect 35897 43775 35955 43781
rect 35897 43741 35909 43775
rect 35943 43741 35955 43775
rect 38562 43772 38568 43784
rect 38523 43744 38568 43772
rect 35897 43735 35955 43741
rect 34480 43676 35204 43704
rect 34480 43664 34486 43676
rect 35526 43664 35532 43716
rect 35584 43664 35590 43716
rect 19705 43639 19763 43645
rect 19705 43605 19717 43639
rect 19751 43636 19763 43639
rect 20622 43636 20628 43648
rect 19751 43608 20628 43636
rect 19751 43605 19763 43608
rect 19705 43599 19763 43605
rect 20622 43596 20628 43608
rect 20680 43636 20686 43648
rect 21174 43636 21180 43648
rect 20680 43608 21180 43636
rect 20680 43596 20686 43608
rect 21174 43596 21180 43608
rect 21232 43596 21238 43648
rect 23014 43636 23020 43648
rect 22975 43608 23020 43636
rect 23014 43596 23020 43608
rect 23072 43596 23078 43648
rect 34606 43596 34612 43648
rect 34664 43636 34670 43648
rect 35912 43636 35940 43735
rect 38562 43732 38568 43744
rect 38620 43732 38626 43784
rect 38654 43732 38660 43784
rect 38712 43772 38718 43784
rect 38712 43744 38757 43772
rect 38712 43732 38718 43744
rect 41138 43636 41144 43648
rect 34664 43608 35940 43636
rect 41099 43608 41144 43636
rect 34664 43596 34670 43608
rect 41138 43596 41144 43608
rect 41196 43596 41202 43648
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 28166 43432 28172 43444
rect 28127 43404 28172 43432
rect 28166 43392 28172 43404
rect 28224 43392 28230 43444
rect 37553 43435 37611 43441
rect 37553 43432 37565 43435
rect 36740 43404 37565 43432
rect 36740 43376 36768 43404
rect 37553 43401 37565 43404
rect 37599 43401 37611 43435
rect 37553 43395 37611 43401
rect 23017 43367 23075 43373
rect 23017 43333 23029 43367
rect 23063 43364 23075 43367
rect 23106 43364 23112 43376
rect 23063 43336 23112 43364
rect 23063 43333 23075 43336
rect 23017 43327 23075 43333
rect 23106 43324 23112 43336
rect 23164 43324 23170 43376
rect 24578 43364 24584 43376
rect 24228 43336 24584 43364
rect 21266 43296 21272 43308
rect 21227 43268 21272 43296
rect 21266 43256 21272 43268
rect 21324 43256 21330 43308
rect 22097 43299 22155 43305
rect 22097 43265 22109 43299
rect 22143 43296 22155 43299
rect 22186 43296 22192 43308
rect 22143 43268 22192 43296
rect 22143 43265 22155 43268
rect 22097 43259 22155 43265
rect 22186 43256 22192 43268
rect 22244 43296 22250 43308
rect 23382 43296 23388 43308
rect 22244 43268 23388 43296
rect 22244 43256 22250 43268
rect 23382 43256 23388 43268
rect 23440 43256 23446 43308
rect 23661 43299 23719 43305
rect 23661 43265 23673 43299
rect 23707 43296 23719 43299
rect 23750 43296 23756 43308
rect 23707 43268 23756 43296
rect 23707 43265 23719 43268
rect 23661 43259 23719 43265
rect 23750 43256 23756 43268
rect 23808 43256 23814 43308
rect 24026 43296 24032 43308
rect 23987 43268 24032 43296
rect 24026 43256 24032 43268
rect 24084 43256 24090 43308
rect 24228 43305 24256 43336
rect 24578 43324 24584 43336
rect 24636 43364 24642 43376
rect 26605 43367 26663 43373
rect 24636 43336 26280 43364
rect 24636 43324 24642 43336
rect 24213 43299 24271 43305
rect 24213 43265 24225 43299
rect 24259 43265 24271 43299
rect 24213 43259 24271 43265
rect 25222 43256 25228 43308
rect 25280 43296 25286 43308
rect 25685 43299 25743 43305
rect 25685 43296 25697 43299
rect 25280 43268 25697 43296
rect 25280 43256 25286 43268
rect 25685 43265 25697 43268
rect 25731 43265 25743 43299
rect 25685 43259 25743 43265
rect 25777 43299 25835 43305
rect 25777 43265 25789 43299
rect 25823 43296 25835 43299
rect 26050 43296 26056 43308
rect 25823 43268 26056 43296
rect 25823 43265 25835 43268
rect 25777 43259 25835 43265
rect 26050 43256 26056 43268
rect 26108 43256 26114 43308
rect 26145 43299 26203 43305
rect 26145 43265 26157 43299
rect 26191 43265 26203 43299
rect 26252 43296 26280 43336
rect 26605 43333 26617 43367
rect 26651 43364 26663 43367
rect 27614 43364 27620 43376
rect 26651 43336 27620 43364
rect 26651 43333 26663 43336
rect 26605 43327 26663 43333
rect 27614 43324 27620 43336
rect 27672 43324 27678 43376
rect 30374 43364 30380 43376
rect 29932 43336 30380 43364
rect 27154 43296 27160 43308
rect 26252 43268 27160 43296
rect 26145 43259 26203 43265
rect 20625 43231 20683 43237
rect 20625 43197 20637 43231
rect 20671 43228 20683 43231
rect 22002 43228 22008 43240
rect 20671 43200 22008 43228
rect 20671 43197 20683 43200
rect 20625 43191 20683 43197
rect 22002 43188 22008 43200
rect 22060 43188 22066 43240
rect 22557 43231 22615 43237
rect 22557 43197 22569 43231
rect 22603 43228 22615 43231
rect 23290 43228 23296 43240
rect 22603 43200 23296 43228
rect 22603 43197 22615 43200
rect 22557 43191 22615 43197
rect 23290 43188 23296 43200
rect 23348 43228 23354 43240
rect 23569 43231 23627 43237
rect 23569 43228 23581 43231
rect 23348 43200 23581 43228
rect 23348 43188 23354 43200
rect 23569 43197 23581 43200
rect 23615 43197 23627 43231
rect 26160 43228 26188 43259
rect 27154 43256 27160 43268
rect 27212 43296 27218 43308
rect 27249 43299 27307 43305
rect 27249 43296 27261 43299
rect 27212 43268 27261 43296
rect 27212 43256 27218 43268
rect 27249 43265 27261 43268
rect 27295 43265 27307 43299
rect 27709 43299 27767 43305
rect 27709 43296 27721 43299
rect 27249 43259 27307 43265
rect 27632 43268 27721 43296
rect 27632 43240 27660 43268
rect 27709 43265 27721 43268
rect 27755 43265 27767 43299
rect 27709 43259 27767 43265
rect 27798 43256 27804 43308
rect 27856 43296 27862 43308
rect 28077 43299 28135 43305
rect 28077 43296 28089 43299
rect 27856 43268 28089 43296
rect 27856 43256 27862 43268
rect 28077 43265 28089 43268
rect 28123 43296 28135 43299
rect 28534 43296 28540 43308
rect 28123 43268 28540 43296
rect 28123 43265 28135 43268
rect 28077 43259 28135 43265
rect 28534 43256 28540 43268
rect 28592 43296 28598 43308
rect 29932 43305 29960 43336
rect 30374 43324 30380 43336
rect 30432 43324 30438 43376
rect 32766 43364 32772 43376
rect 32727 43336 32772 43364
rect 32766 43324 32772 43336
rect 32824 43324 32830 43376
rect 34146 43364 34152 43376
rect 33612 43336 34152 43364
rect 29917 43299 29975 43305
rect 28592 43268 29316 43296
rect 28592 43256 28598 43268
rect 26160 43200 27292 43228
rect 23569 43191 23627 43197
rect 27264 43172 27292 43200
rect 27614 43188 27620 43240
rect 27672 43188 27678 43240
rect 27982 43188 27988 43240
rect 28040 43228 28046 43240
rect 29181 43231 29239 43237
rect 29181 43228 29193 43231
rect 28040 43200 29193 43228
rect 28040 43188 28046 43200
rect 29181 43197 29193 43200
rect 29227 43197 29239 43231
rect 29181 43191 29239 43197
rect 23658 43120 23664 43172
rect 23716 43160 23722 43172
rect 24673 43163 24731 43169
rect 24673 43160 24685 43163
rect 23716 43132 24685 43160
rect 23716 43120 23722 43132
rect 24673 43129 24685 43132
rect 24719 43129 24731 43163
rect 24673 43123 24731 43129
rect 27246 43120 27252 43172
rect 27304 43120 27310 43172
rect 29288 43160 29316 43268
rect 29917 43265 29929 43299
rect 29963 43265 29975 43299
rect 29917 43259 29975 43265
rect 30006 43256 30012 43308
rect 30064 43296 30070 43308
rect 30193 43299 30251 43305
rect 30064 43268 30109 43296
rect 30064 43256 30070 43268
rect 30193 43265 30205 43299
rect 30239 43296 30251 43299
rect 30558 43296 30564 43308
rect 30239 43268 30564 43296
rect 30239 43265 30251 43268
rect 30193 43259 30251 43265
rect 30558 43256 30564 43268
rect 30616 43256 30622 43308
rect 33612 43305 33640 43336
rect 34146 43324 34152 43336
rect 34204 43324 34210 43376
rect 36722 43364 36728 43376
rect 36372 43336 36728 43364
rect 33229 43299 33287 43305
rect 33229 43265 33241 43299
rect 33275 43265 33287 43299
rect 33229 43259 33287 43265
rect 33597 43299 33655 43305
rect 33597 43265 33609 43299
rect 33643 43265 33655 43299
rect 34238 43296 34244 43308
rect 34199 43268 34244 43296
rect 33597 43259 33655 43265
rect 29730 43228 29736 43240
rect 29691 43200 29736 43228
rect 29730 43188 29736 43200
rect 29788 43188 29794 43240
rect 30024 43228 30052 43256
rect 31389 43231 31447 43237
rect 31389 43228 31401 43231
rect 30024 43200 31401 43228
rect 31389 43197 31401 43200
rect 31435 43197 31447 43231
rect 31389 43191 31447 43197
rect 30837 43163 30895 43169
rect 30837 43160 30849 43163
rect 29288 43132 30849 43160
rect 30837 43129 30849 43132
rect 30883 43160 30895 43163
rect 31294 43160 31300 43172
rect 30883 43132 31300 43160
rect 30883 43129 30895 43132
rect 30837 43123 30895 43129
rect 31294 43120 31300 43132
rect 31352 43120 31358 43172
rect 33244 43160 33272 43259
rect 34238 43256 34244 43268
rect 34296 43256 34302 43308
rect 36372 43305 36400 43336
rect 36722 43324 36728 43336
rect 36780 43324 36786 43376
rect 37458 43324 37464 43376
rect 37516 43364 37522 43376
rect 38289 43367 38347 43373
rect 38289 43364 38301 43367
rect 37516 43336 38301 43364
rect 37516 43324 37522 43336
rect 38289 43333 38301 43336
rect 38335 43333 38347 43367
rect 38289 43327 38347 43333
rect 36357 43299 36415 43305
rect 36357 43265 36369 43299
rect 36403 43265 36415 43299
rect 36357 43259 36415 43265
rect 36446 43256 36452 43308
rect 36504 43296 36510 43308
rect 36633 43299 36691 43305
rect 36633 43296 36645 43299
rect 36504 43268 36645 43296
rect 36504 43256 36510 43268
rect 36633 43265 36645 43268
rect 36679 43265 36691 43299
rect 39390 43296 39396 43308
rect 39351 43268 39396 43296
rect 36633 43259 36691 43265
rect 39390 43256 39396 43268
rect 39448 43256 39454 43308
rect 39942 43296 39948 43308
rect 39903 43268 39948 43296
rect 39942 43256 39948 43268
rect 40000 43256 40006 43308
rect 33689 43231 33747 43237
rect 33689 43197 33701 43231
rect 33735 43228 33747 43231
rect 34514 43228 34520 43240
rect 33735 43200 34520 43228
rect 33735 43197 33747 43200
rect 33689 43191 33747 43197
rect 34514 43188 34520 43200
rect 34572 43188 34578 43240
rect 33778 43160 33784 43172
rect 33244 43132 33784 43160
rect 33778 43120 33784 43132
rect 33836 43120 33842 43172
rect 34606 43052 34612 43104
rect 34664 43092 34670 43104
rect 34977 43095 35035 43101
rect 34977 43092 34989 43095
rect 34664 43064 34989 43092
rect 34664 43052 34670 43064
rect 34977 43061 34989 43064
rect 35023 43061 35035 43095
rect 34977 43055 35035 43061
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 23198 42888 23204 42900
rect 23159 42860 23204 42888
rect 23198 42848 23204 42860
rect 23256 42848 23262 42900
rect 25222 42848 25228 42900
rect 25280 42888 25286 42900
rect 25961 42891 26019 42897
rect 25961 42888 25973 42891
rect 25280 42860 25973 42888
rect 25280 42848 25286 42860
rect 22646 42684 22652 42696
rect 22607 42656 22652 42684
rect 22646 42644 22652 42656
rect 22704 42644 22710 42696
rect 23014 42684 23020 42696
rect 22975 42656 23020 42684
rect 23014 42644 23020 42656
rect 23072 42644 23078 42696
rect 25406 42684 25412 42696
rect 25367 42656 25412 42684
rect 25406 42644 25412 42656
rect 25464 42644 25470 42696
rect 25516 42693 25544 42860
rect 25961 42857 25973 42860
rect 26007 42888 26019 42891
rect 26234 42888 26240 42900
rect 26007 42860 26240 42888
rect 26007 42857 26019 42860
rect 25961 42851 26019 42857
rect 26234 42848 26240 42860
rect 26292 42848 26298 42900
rect 29638 42780 29644 42832
rect 29696 42820 29702 42832
rect 30006 42820 30012 42832
rect 29696 42792 30012 42820
rect 29696 42780 29702 42792
rect 30006 42780 30012 42792
rect 30064 42820 30070 42832
rect 31205 42823 31263 42829
rect 31205 42820 31217 42823
rect 30064 42792 31217 42820
rect 30064 42780 30070 42792
rect 27433 42755 27491 42761
rect 27433 42721 27445 42755
rect 27479 42752 27491 42755
rect 28074 42752 28080 42764
rect 27479 42724 28080 42752
rect 27479 42721 27491 42724
rect 27433 42715 27491 42721
rect 28074 42712 28080 42724
rect 28132 42712 28138 42764
rect 28997 42755 29055 42761
rect 28997 42721 29009 42755
rect 29043 42752 29055 42755
rect 29730 42752 29736 42764
rect 29043 42724 29736 42752
rect 29043 42721 29055 42724
rect 28997 42715 29055 42721
rect 29730 42712 29736 42724
rect 29788 42752 29794 42764
rect 30760 42761 30788 42792
rect 31205 42789 31217 42792
rect 31251 42789 31263 42823
rect 31205 42783 31263 42789
rect 30285 42755 30343 42761
rect 30285 42752 30297 42755
rect 29788 42724 30297 42752
rect 29788 42712 29794 42724
rect 30285 42721 30297 42724
rect 30331 42721 30343 42755
rect 30285 42715 30343 42721
rect 30745 42755 30803 42761
rect 30745 42721 30757 42755
rect 30791 42721 30803 42755
rect 33134 42752 33140 42764
rect 33095 42724 33140 42752
rect 30745 42715 30803 42721
rect 33134 42712 33140 42724
rect 33192 42712 33198 42764
rect 33778 42752 33784 42764
rect 33739 42724 33784 42752
rect 33778 42712 33784 42724
rect 33836 42712 33842 42764
rect 34606 42752 34612 42764
rect 34256 42724 34612 42752
rect 25501 42687 25559 42693
rect 25501 42653 25513 42687
rect 25547 42653 25559 42687
rect 25501 42647 25559 42653
rect 27065 42687 27123 42693
rect 27065 42653 27077 42687
rect 27111 42684 27123 42687
rect 27614 42684 27620 42696
rect 27111 42656 27620 42684
rect 27111 42653 27123 42656
rect 27065 42647 27123 42653
rect 27614 42644 27620 42656
rect 27672 42644 27678 42696
rect 27982 42684 27988 42696
rect 27943 42656 27988 42684
rect 27982 42644 27988 42656
rect 28040 42644 28046 42696
rect 28166 42644 28172 42696
rect 28224 42684 28230 42696
rect 28537 42687 28595 42693
rect 28537 42684 28549 42687
rect 28224 42656 28549 42684
rect 28224 42644 28230 42656
rect 28537 42653 28549 42656
rect 28583 42684 28595 42687
rect 28583 42656 28994 42684
rect 28583 42653 28595 42656
rect 28537 42647 28595 42653
rect 23750 42576 23756 42628
rect 23808 42616 23814 42628
rect 24949 42619 25007 42625
rect 24949 42616 24961 42619
rect 23808 42588 24961 42616
rect 23808 42576 23814 42588
rect 24949 42585 24961 42588
rect 24995 42585 25007 42619
rect 24949 42579 25007 42585
rect 26881 42619 26939 42625
rect 26881 42585 26893 42619
rect 26927 42616 26939 42619
rect 27154 42616 27160 42628
rect 26927 42588 27160 42616
rect 26927 42585 26939 42588
rect 26881 42579 26939 42585
rect 27154 42576 27160 42588
rect 27212 42576 27218 42628
rect 22922 42508 22928 42560
rect 22980 42548 22986 42560
rect 28077 42551 28135 42557
rect 28077 42548 28089 42551
rect 22980 42520 28089 42548
rect 22980 42508 22986 42520
rect 28077 42517 28089 42520
rect 28123 42517 28135 42551
rect 28966 42548 28994 42656
rect 30374 42644 30380 42696
rect 30432 42684 30438 42696
rect 30561 42687 30619 42693
rect 30561 42684 30573 42687
rect 30432 42656 30573 42684
rect 30432 42644 30438 42656
rect 30561 42653 30573 42656
rect 30607 42653 30619 42687
rect 32398 42684 32404 42696
rect 32311 42656 32404 42684
rect 30561 42647 30619 42653
rect 32398 42644 32404 42656
rect 32456 42684 32462 42696
rect 33410 42684 33416 42696
rect 32456 42656 33416 42684
rect 32456 42644 32462 42656
rect 33410 42644 33416 42656
rect 33468 42644 33474 42696
rect 34256 42693 34284 42724
rect 34606 42712 34612 42724
rect 34664 42712 34670 42764
rect 34698 42712 34704 42764
rect 34756 42752 34762 42764
rect 34885 42755 34943 42761
rect 34885 42752 34897 42755
rect 34756 42724 34897 42752
rect 34756 42712 34762 42724
rect 34885 42721 34897 42724
rect 34931 42721 34943 42755
rect 34885 42715 34943 42721
rect 35434 42712 35440 42764
rect 35492 42752 35498 42764
rect 35529 42755 35587 42761
rect 35529 42752 35541 42755
rect 35492 42724 35541 42752
rect 35492 42712 35498 42724
rect 35529 42721 35541 42724
rect 35575 42721 35587 42755
rect 35529 42715 35587 42721
rect 36449 42755 36507 42761
rect 36449 42721 36461 42755
rect 36495 42752 36507 42755
rect 37550 42752 37556 42764
rect 36495 42724 37556 42752
rect 36495 42721 36507 42724
rect 36449 42715 36507 42721
rect 37550 42712 37556 42724
rect 37608 42752 37614 42764
rect 38013 42755 38071 42761
rect 38013 42752 38025 42755
rect 37608 42724 38025 42752
rect 37608 42712 37614 42724
rect 38013 42721 38025 42724
rect 38059 42752 38071 42755
rect 38565 42755 38623 42761
rect 38565 42752 38577 42755
rect 38059 42724 38577 42752
rect 38059 42721 38071 42724
rect 38013 42715 38071 42721
rect 38565 42721 38577 42724
rect 38611 42721 38623 42755
rect 38565 42715 38623 42721
rect 39209 42755 39267 42761
rect 39209 42721 39221 42755
rect 39255 42752 39267 42755
rect 40126 42752 40132 42764
rect 39255 42724 40132 42752
rect 39255 42721 39267 42724
rect 39209 42715 39267 42721
rect 40126 42712 40132 42724
rect 40184 42752 40190 42764
rect 41138 42752 41144 42764
rect 40184 42724 41144 42752
rect 40184 42712 40190 42724
rect 41138 42712 41144 42724
rect 41196 42712 41202 42764
rect 34241 42687 34299 42693
rect 34241 42653 34253 42687
rect 34287 42653 34299 42687
rect 34241 42647 34299 42653
rect 34330 42644 34336 42696
rect 34388 42684 34394 42696
rect 34388 42656 34433 42684
rect 34388 42644 34394 42656
rect 37182 42644 37188 42696
rect 37240 42684 37246 42696
rect 37461 42687 37519 42693
rect 37461 42684 37473 42687
rect 37240 42656 37473 42684
rect 37240 42644 37246 42656
rect 37461 42653 37473 42656
rect 37507 42653 37519 42687
rect 37461 42647 37519 42653
rect 29454 42576 29460 42628
rect 29512 42616 29518 42628
rect 29733 42619 29791 42625
rect 29733 42616 29745 42619
rect 29512 42588 29745 42616
rect 29512 42576 29518 42588
rect 29733 42585 29745 42588
rect 29779 42585 29791 42619
rect 29733 42579 29791 42585
rect 30190 42576 30196 42628
rect 30248 42616 30254 42628
rect 30248 42588 30788 42616
rect 30248 42576 30254 42588
rect 30650 42548 30656 42560
rect 28966 42520 30656 42548
rect 28077 42511 28135 42517
rect 30650 42508 30656 42520
rect 30708 42508 30714 42560
rect 30760 42548 30788 42588
rect 31757 42551 31815 42557
rect 31757 42548 31769 42551
rect 30760 42520 31769 42548
rect 31757 42517 31769 42520
rect 31803 42517 31815 42551
rect 36906 42548 36912 42560
rect 36867 42520 36912 42548
rect 31757 42511 31815 42517
rect 36906 42508 36912 42520
rect 36964 42508 36970 42560
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 22646 42304 22652 42356
rect 22704 42344 22710 42356
rect 23661 42347 23719 42353
rect 23661 42344 23673 42347
rect 22704 42316 23673 42344
rect 22704 42304 22710 42316
rect 23661 42313 23673 42316
rect 23707 42313 23719 42347
rect 26234 42344 26240 42356
rect 23661 42307 23719 42313
rect 25332 42316 26240 42344
rect 23750 42208 23756 42220
rect 23711 42180 23756 42208
rect 23750 42168 23756 42180
rect 23808 42168 23814 42220
rect 24026 42168 24032 42220
rect 24084 42208 24090 42220
rect 24305 42211 24363 42217
rect 24305 42208 24317 42211
rect 24084 42180 24317 42208
rect 24084 42168 24090 42180
rect 24305 42177 24317 42180
rect 24351 42208 24363 42211
rect 25133 42211 25191 42217
rect 25133 42208 25145 42211
rect 24351 42180 25145 42208
rect 24351 42177 24363 42180
rect 24305 42171 24363 42177
rect 25133 42177 25145 42180
rect 25179 42177 25191 42211
rect 25332 42208 25360 42316
rect 26234 42304 26240 42316
rect 26292 42304 26298 42356
rect 30101 42347 30159 42353
rect 30101 42344 30113 42347
rect 29104 42316 30113 42344
rect 25406 42236 25412 42288
rect 25464 42276 25470 42288
rect 25464 42248 25728 42276
rect 25464 42236 25470 42248
rect 25700 42217 25728 42248
rect 29104 42217 29132 42316
rect 30101 42313 30113 42316
rect 30147 42344 30159 42347
rect 30558 42344 30564 42356
rect 30147 42316 30564 42344
rect 30147 42313 30159 42316
rect 30101 42307 30159 42313
rect 30558 42304 30564 42316
rect 30616 42304 30622 42356
rect 30650 42304 30656 42356
rect 30708 42344 30714 42356
rect 30708 42316 30753 42344
rect 30708 42304 30714 42316
rect 31018 42304 31024 42356
rect 31076 42344 31082 42356
rect 31757 42347 31815 42353
rect 31757 42344 31769 42347
rect 31076 42316 31769 42344
rect 31076 42304 31082 42316
rect 31757 42313 31769 42316
rect 31803 42344 31815 42347
rect 32309 42347 32367 42353
rect 32309 42344 32321 42347
rect 31803 42316 32321 42344
rect 31803 42313 31815 42316
rect 31757 42307 31815 42313
rect 32309 42313 32321 42316
rect 32355 42313 32367 42347
rect 32309 42307 32367 42313
rect 33873 42347 33931 42353
rect 33873 42313 33885 42347
rect 33919 42344 33931 42347
rect 33962 42344 33968 42356
rect 33919 42316 33968 42344
rect 33919 42313 33931 42316
rect 33873 42307 33931 42313
rect 33962 42304 33968 42316
rect 34020 42304 34026 42356
rect 34330 42304 34336 42356
rect 34388 42344 34394 42356
rect 34425 42347 34483 42353
rect 34425 42344 34437 42347
rect 34388 42316 34437 42344
rect 34388 42304 34394 42316
rect 34425 42313 34437 42316
rect 34471 42344 34483 42347
rect 34977 42347 35035 42353
rect 34977 42344 34989 42347
rect 34471 42316 34989 42344
rect 34471 42313 34483 42316
rect 34425 42307 34483 42313
rect 34977 42313 34989 42316
rect 35023 42344 35035 42347
rect 36173 42347 36231 42353
rect 36173 42344 36185 42347
rect 35023 42316 36185 42344
rect 35023 42313 35035 42316
rect 34977 42307 35035 42313
rect 36173 42313 36185 42316
rect 36219 42344 36231 42347
rect 36906 42344 36912 42356
rect 36219 42316 36912 42344
rect 36219 42313 36231 42316
rect 36173 42307 36231 42313
rect 36906 42304 36912 42316
rect 36964 42304 36970 42356
rect 38102 42344 38108 42356
rect 38063 42316 38108 42344
rect 38102 42304 38108 42316
rect 38160 42304 38166 42356
rect 30576 42276 30604 42304
rect 31113 42279 31171 42285
rect 31113 42276 31125 42279
rect 30576 42248 31125 42276
rect 31113 42245 31125 42248
rect 31159 42245 31171 42279
rect 31113 42239 31171 42245
rect 33321 42279 33379 42285
rect 33321 42245 33333 42279
rect 33367 42276 33379 42279
rect 34348 42276 34376 42304
rect 36722 42276 36728 42288
rect 33367 42248 34376 42276
rect 36683 42248 36728 42276
rect 33367 42245 33379 42248
rect 33321 42239 33379 42245
rect 36722 42236 36728 42248
rect 36780 42276 36786 42288
rect 37461 42279 37519 42285
rect 37461 42276 37473 42279
rect 36780 42248 37473 42276
rect 36780 42236 36786 42248
rect 37461 42245 37473 42248
rect 37507 42245 37519 42279
rect 37461 42239 37519 42245
rect 25501 42211 25559 42217
rect 25501 42208 25513 42211
rect 25332 42180 25513 42208
rect 25133 42171 25191 42177
rect 25501 42177 25513 42180
rect 25547 42177 25559 42211
rect 25501 42171 25559 42177
rect 25685 42211 25743 42217
rect 25685 42177 25697 42211
rect 25731 42208 25743 42211
rect 29089 42211 29147 42217
rect 25731 42180 26648 42208
rect 25731 42177 25743 42180
rect 25685 42171 25743 42177
rect 24578 42140 24584 42152
rect 24539 42112 24584 42140
rect 24578 42100 24584 42112
rect 24636 42100 24642 42152
rect 26620 42016 26648 42180
rect 29089 42177 29101 42211
rect 29135 42177 29147 42211
rect 29454 42208 29460 42220
rect 29415 42180 29460 42208
rect 29089 42171 29147 42177
rect 29454 42168 29460 42180
rect 29512 42168 29518 42220
rect 30650 42168 30656 42220
rect 30708 42208 30714 42220
rect 32214 42208 32220 42220
rect 30708 42180 32220 42208
rect 30708 42168 30714 42180
rect 32214 42168 32220 42180
rect 32272 42168 32278 42220
rect 22002 41964 22008 42016
rect 22060 42004 22066 42016
rect 22649 42007 22707 42013
rect 22649 42004 22661 42007
rect 22060 41976 22661 42004
rect 22060 41964 22066 41976
rect 22649 41973 22661 41976
rect 22695 42004 22707 42007
rect 22738 42004 22744 42016
rect 22695 41976 22744 42004
rect 22695 41973 22707 41976
rect 22649 41967 22707 41973
rect 22738 41964 22744 41976
rect 22796 41964 22802 42016
rect 26602 41964 26608 42016
rect 26660 42004 26666 42016
rect 27617 42007 27675 42013
rect 27617 42004 27629 42007
rect 26660 41976 27629 42004
rect 26660 41964 26666 41976
rect 27617 41973 27629 41976
rect 27663 41973 27675 42007
rect 35526 42004 35532 42016
rect 35487 41976 35532 42004
rect 27617 41967 27675 41973
rect 35526 41964 35532 41976
rect 35584 42004 35590 42016
rect 37182 42004 37188 42016
rect 35584 41976 37188 42004
rect 35584 41964 35590 41976
rect 37182 41964 37188 41976
rect 37240 41964 37246 42016
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 24762 41760 24768 41812
rect 24820 41800 24826 41812
rect 25041 41803 25099 41809
rect 25041 41800 25053 41803
rect 24820 41772 25053 41800
rect 24820 41760 24826 41772
rect 25041 41769 25053 41772
rect 25087 41800 25099 41803
rect 28166 41800 28172 41812
rect 25087 41772 28172 41800
rect 25087 41769 25099 41772
rect 25041 41763 25099 41769
rect 28166 41760 28172 41772
rect 28224 41760 28230 41812
rect 31294 41800 31300 41812
rect 31255 41772 31300 41800
rect 31294 41760 31300 41772
rect 31352 41760 31358 41812
rect 33962 41760 33968 41812
rect 34020 41800 34026 41812
rect 34149 41803 34207 41809
rect 34149 41800 34161 41803
rect 34020 41772 34161 41800
rect 34020 41760 34026 41772
rect 34149 41769 34161 41772
rect 34195 41769 34207 41803
rect 34149 41763 34207 41769
rect 33134 41692 33140 41744
rect 33192 41732 33198 41744
rect 34885 41735 34943 41741
rect 34885 41732 34897 41735
rect 33192 41704 34897 41732
rect 33192 41692 33198 41704
rect 34885 41701 34897 41704
rect 34931 41732 34943 41735
rect 35526 41732 35532 41744
rect 34931 41704 35532 41732
rect 34931 41701 34943 41704
rect 34885 41695 34943 41701
rect 35526 41692 35532 41704
rect 35584 41692 35590 41744
rect 28905 41667 28963 41673
rect 28905 41633 28917 41667
rect 28951 41664 28963 41667
rect 29825 41667 29883 41673
rect 29825 41664 29837 41667
rect 28951 41636 29837 41664
rect 28951 41633 28963 41636
rect 28905 41627 28963 41633
rect 29825 41633 29837 41636
rect 29871 41633 29883 41667
rect 29825 41627 29883 41633
rect 26145 41599 26203 41605
rect 26145 41565 26157 41599
rect 26191 41596 26203 41599
rect 26234 41596 26240 41608
rect 26191 41568 26240 41596
rect 26191 41565 26203 41568
rect 26145 41559 26203 41565
rect 26234 41556 26240 41568
rect 26292 41556 26298 41608
rect 26602 41596 26608 41608
rect 26563 41568 26608 41596
rect 26602 41556 26608 41568
rect 26660 41556 26666 41608
rect 26252 41460 26280 41556
rect 27614 41528 27620 41540
rect 27278 41500 27620 41528
rect 27614 41488 27620 41500
rect 27672 41488 27678 41540
rect 29917 41531 29975 41537
rect 29917 41497 29929 41531
rect 29963 41528 29975 41531
rect 30466 41528 30472 41540
rect 29963 41500 30472 41528
rect 29963 41497 29975 41500
rect 29917 41491 29975 41497
rect 30466 41488 30472 41500
rect 30524 41488 30530 41540
rect 30834 41528 30840 41540
rect 30795 41500 30840 41528
rect 30834 41488 30840 41500
rect 30892 41488 30898 41540
rect 27338 41460 27344 41472
rect 26252 41432 27344 41460
rect 27338 41420 27344 41432
rect 27396 41460 27402 41472
rect 28077 41463 28135 41469
rect 28077 41460 28089 41463
rect 27396 41432 28089 41460
rect 27396 41420 27402 41432
rect 28077 41429 28089 41432
rect 28123 41429 28135 41463
rect 28077 41423 28135 41429
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 22738 41216 22744 41268
rect 22796 41256 22802 41268
rect 24857 41259 24915 41265
rect 24857 41256 24869 41259
rect 22796 41228 24869 41256
rect 22796 41216 22802 41228
rect 24857 41225 24869 41228
rect 24903 41225 24915 41259
rect 24857 41219 24915 41225
rect 26234 41216 26240 41268
rect 26292 41256 26298 41268
rect 26510 41256 26516 41268
rect 26292 41228 26516 41256
rect 26292 41216 26298 41228
rect 26510 41216 26516 41228
rect 26568 41216 26574 41268
rect 27249 41259 27307 41265
rect 27249 41225 27261 41259
rect 27295 41256 27307 41259
rect 27338 41256 27344 41268
rect 27295 41228 27344 41256
rect 27295 41225 27307 41228
rect 27249 41219 27307 41225
rect 27338 41216 27344 41228
rect 27396 41216 27402 41268
rect 28534 41256 28540 41268
rect 28495 41228 28540 41256
rect 28534 41216 28540 41228
rect 28592 41216 28598 41268
rect 29181 41259 29239 41265
rect 29181 41225 29193 41259
rect 29227 41256 29239 41259
rect 32398 41256 32404 41268
rect 29227 41228 32404 41256
rect 29227 41225 29239 41228
rect 29181 41219 29239 41225
rect 32398 41216 32404 41228
rect 32456 41216 32462 41268
rect 25501 41191 25559 41197
rect 25501 41157 25513 41191
rect 25547 41188 25559 41191
rect 25958 41188 25964 41200
rect 25547 41160 25964 41188
rect 25547 41157 25559 41160
rect 25501 41151 25559 41157
rect 25958 41148 25964 41160
rect 26016 41188 26022 41200
rect 27709 41191 27767 41197
rect 27709 41188 27721 41191
rect 26016 41160 27721 41188
rect 26016 41148 26022 41160
rect 27709 41157 27721 41160
rect 27755 41188 27767 41191
rect 30190 41188 30196 41200
rect 27755 41160 30196 41188
rect 27755 41157 27767 41160
rect 27709 41151 27767 41157
rect 30190 41148 30196 41160
rect 30248 41148 30254 41200
rect 26053 41123 26111 41129
rect 26053 41089 26065 41123
rect 26099 41120 26111 41123
rect 26234 41120 26240 41132
rect 26099 41092 26240 41120
rect 26099 41089 26111 41092
rect 26053 41083 26111 41089
rect 26234 41080 26240 41092
rect 26292 41080 26298 41132
rect 29638 40916 29644 40928
rect 29599 40888 29644 40916
rect 29638 40876 29644 40888
rect 29696 40876 29702 40928
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 28813 40715 28871 40721
rect 28813 40681 28825 40715
rect 28859 40712 28871 40715
rect 29638 40712 29644 40724
rect 28859 40684 29644 40712
rect 28859 40681 28871 40684
rect 28813 40675 28871 40681
rect 29638 40672 29644 40684
rect 29696 40672 29702 40724
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 22925 7871 22983 7877
rect 22925 7837 22937 7871
rect 22971 7868 22983 7871
rect 23014 7868 23020 7880
rect 22971 7840 23020 7868
rect 22971 7837 22983 7840
rect 22925 7831 22983 7837
rect 23014 7828 23020 7840
rect 23072 7828 23078 7880
rect 24026 7868 24032 7880
rect 23987 7840 24032 7868
rect 24026 7828 24032 7840
rect 24084 7828 24090 7880
rect 24765 7871 24823 7877
rect 24765 7837 24777 7871
rect 24811 7868 24823 7871
rect 24946 7868 24952 7880
rect 24811 7840 24952 7868
rect 24811 7837 24823 7840
rect 24765 7831 24823 7837
rect 24946 7828 24952 7840
rect 25004 7828 25010 7880
rect 25593 7871 25651 7877
rect 25593 7837 25605 7871
rect 25639 7837 25651 7871
rect 26050 7868 26056 7880
rect 26011 7840 26056 7868
rect 25593 7831 25651 7837
rect 25608 7800 25636 7831
rect 26050 7828 26056 7840
rect 26108 7828 26114 7880
rect 26142 7800 26148 7812
rect 25608 7772 26148 7800
rect 26142 7760 26148 7772
rect 26200 7760 26206 7812
rect 25406 7732 25412 7744
rect 25367 7704 25412 7732
rect 25406 7692 25412 7704
rect 25464 7692 25470 7744
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 21266 7528 21272 7540
rect 21227 7500 21272 7528
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 24854 7460 24860 7472
rect 24815 7432 24860 7460
rect 24854 7420 24860 7432
rect 24912 7420 24918 7472
rect 24946 7420 24952 7472
rect 25004 7460 25010 7472
rect 25682 7460 25688 7472
rect 25004 7432 25049 7460
rect 25643 7432 25688 7460
rect 25004 7420 25010 7432
rect 25682 7420 25688 7432
rect 25740 7420 25746 7472
rect 22094 7352 22100 7404
rect 22152 7392 22158 7404
rect 22649 7395 22707 7401
rect 22649 7392 22661 7395
rect 22152 7364 22661 7392
rect 22152 7352 22158 7364
rect 22649 7361 22661 7364
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 24673 7327 24731 7333
rect 24673 7293 24685 7327
rect 24719 7324 24731 7327
rect 25222 7324 25228 7336
rect 24719 7296 25228 7324
rect 24719 7293 24731 7296
rect 24673 7287 24731 7293
rect 25222 7284 25228 7296
rect 25280 7284 25286 7336
rect 25593 7327 25651 7333
rect 25593 7293 25605 7327
rect 25639 7324 25651 7327
rect 26050 7324 26056 7336
rect 25639 7296 26056 7324
rect 25639 7293 25651 7296
rect 25593 7287 25651 7293
rect 26050 7284 26056 7296
rect 26108 7284 26114 7336
rect 26602 7324 26608 7336
rect 26563 7296 26608 7324
rect 26602 7284 26608 7296
rect 26660 7284 26666 7336
rect 22189 7191 22247 7197
rect 22189 7157 22201 7191
rect 22235 7188 22247 7191
rect 22462 7188 22468 7200
rect 22235 7160 22468 7188
rect 22235 7157 22247 7160
rect 22189 7151 22247 7157
rect 22462 7148 22468 7160
rect 22520 7148 22526 7200
rect 22925 7191 22983 7197
rect 22925 7157 22937 7191
rect 22971 7188 22983 7191
rect 23106 7188 23112 7200
rect 22971 7160 23112 7188
rect 22971 7157 22983 7160
rect 22925 7151 22983 7157
rect 23106 7148 23112 7160
rect 23164 7148 23170 7200
rect 26234 7148 26240 7200
rect 26292 7188 26298 7200
rect 27157 7191 27215 7197
rect 27157 7188 27169 7191
rect 26292 7160 27169 7188
rect 26292 7148 26298 7160
rect 27157 7157 27169 7160
rect 27203 7157 27215 7191
rect 27157 7151 27215 7157
rect 27706 7148 27712 7200
rect 27764 7188 27770 7200
rect 27801 7191 27859 7197
rect 27801 7188 27813 7191
rect 27764 7160 27813 7188
rect 27764 7148 27770 7160
rect 27801 7157 27813 7160
rect 27847 7157 27859 7191
rect 27801 7151 27859 7157
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 24854 6984 24860 6996
rect 24815 6956 24860 6984
rect 24854 6944 24860 6956
rect 24912 6944 24918 6996
rect 25682 6984 25688 6996
rect 25643 6956 25688 6984
rect 25682 6944 25688 6956
rect 25740 6944 25746 6996
rect 23014 6848 23020 6860
rect 22975 6820 23020 6848
rect 23014 6808 23020 6820
rect 23072 6808 23078 6860
rect 23842 6848 23848 6860
rect 23803 6820 23848 6848
rect 23842 6808 23848 6820
rect 23900 6808 23906 6860
rect 27706 6848 27712 6860
rect 27667 6820 27712 6848
rect 27706 6808 27712 6820
rect 27764 6808 27770 6860
rect 27982 6848 27988 6860
rect 27943 6820 27988 6848
rect 27982 6808 27988 6820
rect 28040 6808 28046 6860
rect 20717 6783 20775 6789
rect 20717 6780 20729 6783
rect 20180 6752 20729 6780
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 20180 6653 20208 6752
rect 20717 6749 20729 6752
rect 20763 6780 20775 6783
rect 21266 6780 21272 6792
rect 20763 6752 21272 6780
rect 20763 6749 20775 6752
rect 20717 6743 20775 6749
rect 21266 6740 21272 6752
rect 21324 6780 21330 6792
rect 21453 6783 21511 6789
rect 21453 6780 21465 6783
rect 21324 6752 21465 6780
rect 21324 6740 21330 6752
rect 21453 6749 21465 6752
rect 21499 6749 21511 6783
rect 21453 6743 21511 6749
rect 22465 6783 22523 6789
rect 22465 6749 22477 6783
rect 22511 6749 22523 6783
rect 22465 6743 22523 6749
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6749 24639 6783
rect 24581 6743 24639 6749
rect 22480 6712 22508 6743
rect 20916 6684 22508 6712
rect 20916 6656 20944 6684
rect 20165 6647 20223 6653
rect 20165 6644 20177 6647
rect 19392 6616 20177 6644
rect 19392 6604 19398 6616
rect 20165 6613 20177 6616
rect 20211 6613 20223 6647
rect 20898 6644 20904 6656
rect 20859 6616 20904 6644
rect 20165 6607 20223 6613
rect 20898 6604 20904 6616
rect 20956 6604 20962 6656
rect 21542 6604 21548 6656
rect 21600 6644 21606 6656
rect 21637 6647 21695 6653
rect 21637 6644 21649 6647
rect 21600 6616 21649 6644
rect 21600 6604 21606 6616
rect 21637 6613 21649 6616
rect 21683 6644 21695 6647
rect 22094 6644 22100 6656
rect 21683 6616 22100 6644
rect 21683 6613 21695 6616
rect 21637 6607 21695 6613
rect 22094 6604 22100 6616
rect 22152 6604 22158 6656
rect 22278 6644 22284 6656
rect 22239 6616 22284 6644
rect 22278 6604 22284 6616
rect 22336 6604 22342 6656
rect 22480 6644 22508 6684
rect 23106 6672 23112 6724
rect 23164 6712 23170 6724
rect 23164 6684 23209 6712
rect 23164 6672 23170 6684
rect 23382 6672 23388 6724
rect 23440 6712 23446 6724
rect 24596 6712 24624 6743
rect 25406 6740 25412 6792
rect 25464 6780 25470 6792
rect 25685 6783 25743 6789
rect 25685 6780 25697 6783
rect 25464 6752 25697 6780
rect 25464 6740 25470 6752
rect 25685 6749 25697 6752
rect 25731 6749 25743 6783
rect 25685 6743 25743 6749
rect 26421 6783 26479 6789
rect 26421 6749 26433 6783
rect 26467 6749 26479 6783
rect 26421 6743 26479 6749
rect 23440 6684 24624 6712
rect 23440 6672 23446 6684
rect 26142 6644 26148 6656
rect 22480 6616 26148 6644
rect 26142 6604 26148 6616
rect 26200 6644 26206 6656
rect 26436 6644 26464 6743
rect 27798 6712 27804 6724
rect 27759 6684 27804 6712
rect 27798 6672 27804 6684
rect 27856 6672 27862 6724
rect 26200 6616 26464 6644
rect 26605 6647 26663 6653
rect 26200 6604 26206 6616
rect 26605 6613 26617 6647
rect 26651 6644 26663 6647
rect 28994 6644 29000 6656
rect 26651 6616 29000 6644
rect 26651 6613 26663 6616
rect 26605 6607 26663 6613
rect 28994 6604 29000 6616
rect 29052 6604 29058 6656
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 27617 6443 27675 6449
rect 27617 6409 27629 6443
rect 27663 6440 27675 6443
rect 27798 6440 27804 6452
rect 27663 6412 27804 6440
rect 27663 6409 27675 6412
rect 27617 6403 27675 6409
rect 27798 6400 27804 6412
rect 27856 6400 27862 6452
rect 20530 6372 20536 6384
rect 20491 6344 20536 6372
rect 20530 6332 20536 6344
rect 20588 6332 20594 6384
rect 22554 6372 22560 6384
rect 22515 6344 22560 6372
rect 22554 6332 22560 6344
rect 22612 6332 22618 6384
rect 24026 6372 24032 6384
rect 23987 6344 24032 6372
rect 24026 6332 24032 6344
rect 24084 6332 24090 6384
rect 24118 6332 24124 6384
rect 24176 6372 24182 6384
rect 25682 6372 25688 6384
rect 24176 6344 24221 6372
rect 25643 6344 25688 6372
rect 24176 6332 24182 6344
rect 25682 6332 25688 6344
rect 25740 6332 25746 6384
rect 26510 6264 26516 6316
rect 26568 6304 26574 6316
rect 27617 6307 27675 6313
rect 27617 6304 27629 6307
rect 26568 6276 27629 6304
rect 26568 6264 26574 6276
rect 27617 6273 27629 6276
rect 27663 6304 27675 6307
rect 28261 6307 28319 6313
rect 28261 6304 28273 6307
rect 27663 6276 28273 6304
rect 27663 6273 27675 6276
rect 27617 6267 27675 6273
rect 28261 6273 28273 6276
rect 28307 6273 28319 6307
rect 28261 6267 28319 6273
rect 19889 6239 19947 6245
rect 19889 6205 19901 6239
rect 19935 6236 19947 6239
rect 20441 6239 20499 6245
rect 20441 6236 20453 6239
rect 19935 6208 20453 6236
rect 19935 6205 19947 6208
rect 19889 6199 19947 6205
rect 20441 6205 20453 6208
rect 20487 6205 20499 6239
rect 21082 6236 21088 6248
rect 21043 6208 21088 6236
rect 20441 6199 20499 6205
rect 21082 6196 21088 6208
rect 21140 6196 21146 6248
rect 22462 6236 22468 6248
rect 22423 6208 22468 6236
rect 22462 6196 22468 6208
rect 22520 6196 22526 6248
rect 23477 6239 23535 6245
rect 23477 6205 23489 6239
rect 23523 6236 23535 6239
rect 23566 6236 23572 6248
rect 23523 6208 23572 6236
rect 23523 6205 23535 6208
rect 23477 6199 23535 6205
rect 23566 6196 23572 6208
rect 23624 6196 23630 6248
rect 24946 6236 24952 6248
rect 24907 6208 24952 6236
rect 24946 6196 24952 6208
rect 25004 6196 25010 6248
rect 25593 6239 25651 6245
rect 25593 6205 25605 6239
rect 25639 6236 25651 6239
rect 26234 6236 26240 6248
rect 25639 6208 26240 6236
rect 25639 6205 25651 6208
rect 25593 6199 25651 6205
rect 26234 6196 26240 6208
rect 26292 6196 26298 6248
rect 26421 6239 26479 6245
rect 26421 6236 26433 6239
rect 26344 6208 26433 6236
rect 26344 6180 26372 6208
rect 26421 6205 26433 6208
rect 26467 6205 26479 6239
rect 26421 6199 26479 6205
rect 26326 6128 26332 6180
rect 26384 6128 26390 6180
rect 28166 6060 28172 6112
rect 28224 6100 28230 6112
rect 28261 6103 28319 6109
rect 28261 6100 28273 6103
rect 28224 6072 28273 6100
rect 28224 6060 28230 6072
rect 28261 6069 28273 6072
rect 28307 6069 28319 6103
rect 28261 6063 28319 6069
rect 29181 6103 29239 6109
rect 29181 6069 29193 6103
rect 29227 6100 29239 6103
rect 29730 6100 29736 6112
rect 29227 6072 29736 6100
rect 29227 6069 29239 6072
rect 29181 6063 29239 6069
rect 29730 6060 29736 6072
rect 29788 6060 29794 6112
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 20530 5856 20536 5908
rect 20588 5896 20594 5908
rect 20809 5899 20867 5905
rect 20809 5896 20821 5899
rect 20588 5868 20821 5896
rect 20588 5856 20594 5868
rect 20809 5865 20821 5868
rect 20855 5865 20867 5899
rect 22554 5896 22560 5908
rect 22515 5868 22560 5896
rect 20809 5859 20867 5865
rect 22554 5856 22560 5868
rect 22612 5856 22618 5908
rect 24118 5856 24124 5908
rect 24176 5896 24182 5908
rect 24673 5899 24731 5905
rect 24673 5896 24685 5899
rect 24176 5868 24685 5896
rect 24176 5856 24182 5868
rect 24673 5865 24685 5868
rect 24719 5865 24731 5899
rect 25682 5896 25688 5908
rect 25643 5868 25688 5896
rect 24673 5859 24731 5865
rect 25682 5856 25688 5868
rect 25740 5856 25746 5908
rect 26421 5899 26479 5905
rect 26421 5865 26433 5899
rect 26467 5896 26479 5899
rect 26510 5896 26516 5908
rect 26467 5868 26516 5896
rect 26467 5865 26479 5868
rect 26421 5859 26479 5865
rect 26510 5856 26516 5868
rect 26568 5856 26574 5908
rect 22278 5720 22284 5772
rect 22336 5760 22342 5772
rect 22336 5732 22876 5760
rect 22336 5720 22342 5732
rect 22848 5704 22876 5732
rect 26142 5720 26148 5772
rect 26200 5760 26206 5772
rect 27706 5760 27712 5772
rect 26200 5732 26280 5760
rect 27667 5732 27712 5760
rect 26200 5720 26206 5732
rect 20165 5695 20223 5701
rect 20165 5661 20177 5695
rect 20211 5692 20223 5695
rect 20346 5692 20352 5704
rect 20211 5664 20352 5692
rect 20211 5661 20223 5664
rect 20165 5655 20223 5661
rect 20346 5652 20352 5664
rect 20404 5652 20410 5704
rect 20898 5692 20904 5704
rect 20859 5664 20904 5692
rect 20898 5652 20904 5664
rect 20956 5652 20962 5704
rect 21542 5652 21548 5704
rect 21600 5692 21606 5704
rect 21637 5695 21695 5701
rect 21637 5692 21649 5695
rect 21600 5664 21649 5692
rect 21600 5652 21606 5664
rect 21637 5661 21649 5664
rect 21683 5692 21695 5695
rect 22557 5695 22615 5701
rect 22557 5692 22569 5695
rect 21683 5664 22569 5692
rect 21683 5661 21695 5664
rect 21637 5655 21695 5661
rect 22557 5661 22569 5664
rect 22603 5661 22615 5695
rect 22557 5655 22615 5661
rect 22830 5652 22836 5704
rect 22888 5692 22894 5704
rect 23382 5692 23388 5704
rect 22888 5664 23388 5692
rect 22888 5652 22894 5664
rect 23382 5652 23388 5664
rect 23440 5692 23446 5704
rect 23661 5695 23719 5701
rect 23661 5692 23673 5695
rect 23440 5664 23673 5692
rect 23440 5652 23446 5664
rect 23661 5661 23673 5664
rect 23707 5692 23719 5695
rect 24673 5695 24731 5701
rect 24673 5692 24685 5695
rect 23707 5664 24685 5692
rect 23707 5661 23719 5664
rect 23661 5655 23719 5661
rect 24673 5661 24685 5664
rect 24719 5661 24731 5695
rect 25406 5692 25412 5704
rect 25367 5664 25412 5692
rect 24673 5655 24731 5661
rect 25406 5652 25412 5664
rect 25464 5652 25470 5704
rect 26252 5701 26280 5732
rect 27706 5720 27712 5732
rect 27764 5720 27770 5772
rect 26237 5695 26295 5701
rect 26237 5661 26249 5695
rect 26283 5661 26295 5695
rect 28994 5692 29000 5704
rect 28955 5664 29000 5692
rect 26237 5655 26295 5661
rect 28994 5652 29000 5664
rect 29052 5652 29058 5704
rect 22005 5627 22063 5633
rect 22005 5593 22017 5627
rect 22051 5624 22063 5627
rect 22646 5624 22652 5636
rect 22051 5596 22652 5624
rect 22051 5593 22063 5596
rect 22005 5587 22063 5593
rect 22646 5584 22652 5596
rect 22704 5584 22710 5636
rect 24029 5627 24087 5633
rect 24029 5593 24041 5627
rect 24075 5624 24087 5627
rect 24302 5624 24308 5636
rect 24075 5596 24308 5624
rect 24075 5593 24087 5596
rect 24029 5587 24087 5593
rect 24302 5584 24308 5596
rect 24360 5584 24366 5636
rect 28166 5624 28172 5636
rect 28127 5596 28172 5624
rect 28166 5584 28172 5596
rect 28224 5584 28230 5636
rect 28258 5584 28264 5636
rect 28316 5624 28322 5636
rect 29181 5627 29239 5633
rect 28316 5596 28361 5624
rect 28316 5584 28322 5596
rect 29181 5593 29193 5627
rect 29227 5624 29239 5627
rect 29638 5624 29644 5636
rect 29227 5596 29644 5624
rect 29227 5593 29239 5596
rect 29181 5587 29239 5593
rect 29638 5584 29644 5596
rect 29696 5584 29702 5636
rect 20070 5556 20076 5568
rect 20031 5528 20076 5556
rect 20070 5516 20076 5528
rect 20128 5516 20134 5568
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 19889 5287 19947 5293
rect 19889 5253 19901 5287
rect 19935 5284 19947 5287
rect 20070 5284 20076 5296
rect 19935 5256 20076 5284
rect 19935 5253 19947 5256
rect 19889 5247 19947 5253
rect 20070 5244 20076 5256
rect 20128 5244 20134 5296
rect 22646 5284 22652 5296
rect 22607 5256 22652 5284
rect 22646 5244 22652 5256
rect 22704 5244 22710 5296
rect 24302 5284 24308 5296
rect 24263 5256 24308 5284
rect 24302 5244 24308 5256
rect 24360 5244 24366 5296
rect 26605 5287 26663 5293
rect 26605 5253 26617 5287
rect 26651 5284 26663 5287
rect 27341 5287 27399 5293
rect 27341 5284 27353 5287
rect 26651 5256 27353 5284
rect 26651 5253 26663 5256
rect 26605 5247 26663 5253
rect 27341 5253 27353 5256
rect 27387 5253 27399 5287
rect 29638 5284 29644 5296
rect 29599 5256 29644 5284
rect 27341 5247 27399 5253
rect 29638 5244 29644 5256
rect 29696 5244 29702 5296
rect 29730 5244 29736 5296
rect 29788 5284 29794 5296
rect 29788 5256 29833 5284
rect 29788 5244 29794 5256
rect 26510 5216 26516 5228
rect 26471 5188 26516 5216
rect 26510 5176 26516 5188
rect 26568 5176 26574 5228
rect 18230 5108 18236 5160
rect 18288 5148 18294 5160
rect 19797 5151 19855 5157
rect 19797 5148 19809 5151
rect 18288 5120 19809 5148
rect 18288 5108 18294 5120
rect 19797 5117 19809 5120
rect 19843 5117 19855 5151
rect 19797 5111 19855 5117
rect 20809 5151 20867 5157
rect 20809 5117 20821 5151
rect 20855 5148 20867 5151
rect 21634 5148 21640 5160
rect 20855 5120 21640 5148
rect 20855 5117 20867 5120
rect 20809 5111 20867 5117
rect 21634 5108 21640 5120
rect 21692 5108 21698 5160
rect 22554 5148 22560 5160
rect 22515 5120 22560 5148
rect 22554 5108 22560 5120
rect 22612 5108 22618 5160
rect 23198 5148 23204 5160
rect 23159 5120 23204 5148
rect 23198 5108 23204 5120
rect 23256 5108 23262 5160
rect 24213 5151 24271 5157
rect 24213 5117 24225 5151
rect 24259 5117 24271 5151
rect 24854 5148 24860 5160
rect 24815 5120 24860 5148
rect 24213 5111 24271 5117
rect 21453 5083 21511 5089
rect 21453 5049 21465 5083
rect 21499 5080 21511 5083
rect 24228 5080 24256 5111
rect 24854 5108 24860 5120
rect 24912 5108 24918 5160
rect 27246 5148 27252 5160
rect 27207 5120 27252 5148
rect 27246 5108 27252 5120
rect 27304 5108 27310 5160
rect 27614 5148 27620 5160
rect 27575 5120 27620 5148
rect 27614 5108 27620 5120
rect 27672 5108 27678 5160
rect 28810 5148 28816 5160
rect 28771 5120 28816 5148
rect 28810 5108 28816 5120
rect 28868 5108 28874 5160
rect 21499 5052 24256 5080
rect 21499 5049 21511 5052
rect 21453 5043 21511 5049
rect 19245 5015 19303 5021
rect 19245 4981 19257 5015
rect 19291 5012 19303 5015
rect 21174 5012 21180 5024
rect 19291 4984 21180 5012
rect 19291 4981 19303 4984
rect 19245 4975 19303 4981
rect 21174 4972 21180 4984
rect 21232 4972 21238 5024
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 18230 4808 18236 4820
rect 18191 4780 18236 4808
rect 18230 4768 18236 4780
rect 18288 4768 18294 4820
rect 18877 4811 18935 4817
rect 18877 4777 18889 4811
rect 18923 4808 18935 4811
rect 22554 4808 22560 4820
rect 18923 4780 22560 4808
rect 18923 4777 18935 4780
rect 18877 4771 18935 4777
rect 22554 4768 22560 4780
rect 22612 4768 22618 4820
rect 24765 4811 24823 4817
rect 24765 4777 24777 4811
rect 24811 4808 24823 4811
rect 27246 4808 27252 4820
rect 24811 4780 27252 4808
rect 24811 4777 24823 4780
rect 24765 4771 24823 4777
rect 27246 4768 27252 4780
rect 27304 4768 27310 4820
rect 27433 4811 27491 4817
rect 27433 4777 27445 4811
rect 27479 4808 27491 4811
rect 28258 4808 28264 4820
rect 27479 4780 28264 4808
rect 27479 4777 27491 4780
rect 27433 4771 27491 4777
rect 28258 4768 28264 4780
rect 28316 4768 28322 4820
rect 21174 4672 21180 4684
rect 21135 4644 21180 4672
rect 21174 4632 21180 4644
rect 21232 4632 21238 4684
rect 21818 4672 21824 4684
rect 21779 4644 21824 4672
rect 21818 4632 21824 4644
rect 21876 4632 21882 4684
rect 25498 4672 25504 4684
rect 23952 4644 25504 4672
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19521 4607 19579 4613
rect 19521 4604 19533 4607
rect 19392 4576 19533 4604
rect 19392 4564 19398 4576
rect 19521 4573 19533 4576
rect 19567 4573 19579 4607
rect 20346 4604 20352 4616
rect 20307 4576 20352 4604
rect 19521 4567 19579 4573
rect 20346 4564 20352 4576
rect 20404 4564 20410 4616
rect 22830 4604 22836 4616
rect 22791 4576 22836 4604
rect 22830 4564 22836 4576
rect 22888 4564 22894 4616
rect 23952 4613 23980 4644
rect 25498 4632 25504 4644
rect 25556 4632 25562 4684
rect 25958 4672 25964 4684
rect 25919 4644 25964 4672
rect 25958 4632 25964 4644
rect 26016 4632 26022 4684
rect 28813 4675 28871 4681
rect 28813 4641 28825 4675
rect 28859 4672 28871 4675
rect 28994 4672 29000 4684
rect 28859 4644 29000 4672
rect 28859 4641 28871 4644
rect 28813 4635 28871 4641
rect 28994 4632 29000 4644
rect 29052 4632 29058 4684
rect 29089 4675 29147 4681
rect 29089 4641 29101 4675
rect 29135 4672 29147 4675
rect 30561 4675 30619 4681
rect 30561 4672 30573 4675
rect 29135 4644 30573 4672
rect 29135 4641 29147 4644
rect 29089 4635 29147 4641
rect 30561 4641 30573 4644
rect 30607 4641 30619 4675
rect 30561 4635 30619 4641
rect 23937 4607 23995 4613
rect 23937 4573 23949 4607
rect 23983 4573 23995 4607
rect 23937 4567 23995 4573
rect 29270 4564 29276 4616
rect 29328 4604 29334 4616
rect 29825 4607 29883 4613
rect 29825 4604 29837 4607
rect 29328 4576 29837 4604
rect 29328 4564 29334 4576
rect 29825 4573 29837 4576
rect 29871 4604 29883 4607
rect 30098 4604 30104 4616
rect 29871 4576 30104 4604
rect 29871 4573 29883 4576
rect 29825 4567 29883 4573
rect 30098 4564 30104 4576
rect 30156 4564 30162 4616
rect 21269 4539 21327 4545
rect 21269 4505 21281 4539
rect 21315 4505 21327 4539
rect 21269 4499 21327 4505
rect 23201 4539 23259 4545
rect 23201 4505 23213 4539
rect 23247 4536 23259 4539
rect 23474 4536 23480 4548
rect 23247 4508 23480 4536
rect 23247 4505 23259 4508
rect 23201 4499 23259 4505
rect 19705 4471 19763 4477
rect 19705 4437 19717 4471
rect 19751 4468 19763 4471
rect 20346 4468 20352 4480
rect 19751 4440 20352 4468
rect 19751 4437 19763 4440
rect 19705 4431 19763 4437
rect 20346 4428 20352 4440
rect 20404 4428 20410 4480
rect 20533 4471 20591 4477
rect 20533 4437 20545 4471
rect 20579 4468 20591 4471
rect 21284 4468 21312 4499
rect 23474 4496 23480 4508
rect 23532 4496 23538 4548
rect 24029 4539 24087 4545
rect 24029 4505 24041 4539
rect 24075 4536 24087 4539
rect 25038 4536 25044 4548
rect 24075 4508 25044 4536
rect 24075 4505 24087 4508
rect 24029 4499 24087 4505
rect 25038 4496 25044 4508
rect 25096 4496 25102 4548
rect 25317 4539 25375 4545
rect 25317 4505 25329 4539
rect 25363 4505 25375 4539
rect 25317 4499 25375 4505
rect 20579 4440 21312 4468
rect 25332 4468 25360 4499
rect 25406 4496 25412 4548
rect 25464 4536 25470 4548
rect 28997 4539 29055 4545
rect 25464 4508 25509 4536
rect 25464 4496 25470 4508
rect 28997 4505 29009 4539
rect 29043 4505 29055 4539
rect 28997 4499 29055 4505
rect 26418 4468 26424 4480
rect 25332 4440 26424 4468
rect 20579 4437 20591 4440
rect 20533 4431 20591 4437
rect 26418 4428 26424 4440
rect 26476 4428 26482 4480
rect 29012 4468 29040 4499
rect 29825 4471 29883 4477
rect 29825 4468 29837 4471
rect 29012 4440 29837 4468
rect 29825 4437 29837 4440
rect 29871 4437 29883 4471
rect 29825 4431 29883 4437
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 22830 4264 22836 4276
rect 21284 4236 22836 4264
rect 20346 4128 20352 4140
rect 20307 4100 20352 4128
rect 20346 4088 20352 4100
rect 20404 4088 20410 4140
rect 21284 4137 21312 4236
rect 22830 4224 22836 4236
rect 22888 4224 22894 4276
rect 25406 4264 25412 4276
rect 25367 4236 25412 4264
rect 25406 4224 25412 4236
rect 25464 4224 25470 4276
rect 22189 4199 22247 4205
rect 22189 4196 22201 4199
rect 21928 4168 22201 4196
rect 21269 4131 21327 4137
rect 21269 4097 21281 4131
rect 21315 4097 21327 4131
rect 21269 4091 21327 4097
rect 21450 4088 21456 4140
rect 21508 4128 21514 4140
rect 21928 4128 21956 4168
rect 22189 4165 22201 4168
rect 22235 4165 22247 4199
rect 22189 4159 22247 4165
rect 23474 4156 23480 4208
rect 23532 4196 23538 4208
rect 23753 4199 23811 4205
rect 23753 4196 23765 4199
rect 23532 4168 23765 4196
rect 23532 4156 23538 4168
rect 23753 4165 23765 4168
rect 23799 4165 23811 4199
rect 28077 4199 28135 4205
rect 28077 4196 28089 4199
rect 23753 4159 23811 4165
rect 27356 4168 28089 4196
rect 25498 4128 25504 4140
rect 21508 4100 21956 4128
rect 25459 4100 25504 4128
rect 21508 4088 21514 4100
rect 25498 4088 25504 4100
rect 25556 4088 25562 4140
rect 26510 4128 26516 4140
rect 26471 4100 26516 4128
rect 26510 4088 26516 4100
rect 26568 4088 26574 4140
rect 26605 4131 26663 4137
rect 26605 4097 26617 4131
rect 26651 4128 26663 4131
rect 27356 4128 27384 4168
rect 28077 4165 28089 4168
rect 28123 4165 28135 4199
rect 28077 4159 28135 4165
rect 26651 4100 27384 4128
rect 29089 4131 29147 4137
rect 26651 4097 26663 4100
rect 26605 4091 26663 4097
rect 29089 4097 29101 4131
rect 29135 4128 29147 4131
rect 29178 4128 29184 4140
rect 29135 4100 29184 4128
rect 29135 4097 29147 4100
rect 29089 4091 29147 4097
rect 29178 4088 29184 4100
rect 29236 4088 29242 4140
rect 19153 4063 19211 4069
rect 19153 4029 19165 4063
rect 19199 4060 19211 4063
rect 22097 4063 22155 4069
rect 22097 4060 22109 4063
rect 19199 4032 22109 4060
rect 19199 4029 19211 4032
rect 19153 4023 19211 4029
rect 22097 4029 22109 4032
rect 22143 4029 22155 4063
rect 22097 4023 22155 4029
rect 22278 4020 22284 4072
rect 22336 4060 22342 4072
rect 22373 4063 22431 4069
rect 22373 4060 22385 4063
rect 22336 4032 22385 4060
rect 22336 4020 22342 4032
rect 22373 4029 22385 4032
rect 22419 4029 22431 4063
rect 22373 4023 22431 4029
rect 23661 4063 23719 4069
rect 23661 4029 23673 4063
rect 23707 4029 23719 4063
rect 24118 4060 24124 4072
rect 24079 4032 24124 4060
rect 23661 4023 23719 4029
rect 17865 3995 17923 4001
rect 17865 3961 17877 3995
rect 17911 3992 17923 3995
rect 18598 3992 18604 4004
rect 17911 3964 18604 3992
rect 17911 3961 17923 3964
rect 17865 3955 17923 3961
rect 18598 3952 18604 3964
rect 18656 3952 18662 4004
rect 19797 3995 19855 4001
rect 19797 3961 19809 3995
rect 19843 3992 19855 3995
rect 23676 3992 23704 4023
rect 24118 4020 24124 4032
rect 24176 4020 24182 4072
rect 26878 4020 26884 4072
rect 26936 4060 26942 4072
rect 27157 4063 27215 4069
rect 27157 4060 27169 4063
rect 26936 4032 27169 4060
rect 26936 4020 26942 4032
rect 27157 4029 27169 4032
rect 27203 4029 27215 4063
rect 27157 4023 27215 4029
rect 28169 4063 28227 4069
rect 28169 4029 28181 4063
rect 28215 4060 28227 4063
rect 29549 4063 29607 4069
rect 29549 4060 29561 4063
rect 28215 4032 29561 4060
rect 28215 4029 28227 4032
rect 28169 4023 28227 4029
rect 29549 4029 29561 4032
rect 29595 4029 29607 4063
rect 29549 4023 29607 4029
rect 19843 3964 23704 3992
rect 19843 3961 19855 3964
rect 19797 3955 19855 3961
rect 16114 3924 16120 3936
rect 16075 3896 16120 3924
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 17218 3924 17224 3936
rect 17179 3896 17224 3924
rect 17218 3884 17224 3896
rect 17276 3884 17282 3936
rect 18509 3927 18567 3933
rect 18509 3893 18521 3927
rect 18555 3924 18567 3927
rect 19426 3924 19432 3936
rect 18555 3896 19432 3924
rect 18555 3893 18567 3896
rect 18509 3887 18567 3893
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 20533 3927 20591 3933
rect 20533 3893 20545 3927
rect 20579 3924 20591 3927
rect 21266 3924 21272 3936
rect 20579 3896 21272 3924
rect 20579 3893 20591 3896
rect 20533 3887 20591 3893
rect 21266 3884 21272 3896
rect 21324 3884 21330 3936
rect 21361 3927 21419 3933
rect 21361 3893 21373 3927
rect 21407 3924 21419 3927
rect 23750 3924 23756 3936
rect 21407 3896 23756 3924
rect 21407 3893 21419 3896
rect 21361 3887 21419 3893
rect 23750 3884 23756 3896
rect 23808 3884 23814 3936
rect 28718 3884 28724 3936
rect 28776 3924 28782 3936
rect 28813 3927 28871 3933
rect 28813 3924 28825 3927
rect 28776 3896 28825 3924
rect 28776 3884 28782 3896
rect 28813 3893 28825 3896
rect 28859 3893 28871 3927
rect 30190 3924 30196 3936
rect 30151 3896 30196 3924
rect 28813 3887 28871 3893
rect 30190 3884 30196 3896
rect 30248 3884 30254 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 18233 3723 18291 3729
rect 18233 3689 18245 3723
rect 18279 3720 18291 3723
rect 20070 3720 20076 3732
rect 18279 3692 20076 3720
rect 18279 3689 18291 3692
rect 18233 3683 18291 3689
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 16301 3655 16359 3661
rect 16301 3621 16313 3655
rect 16347 3652 16359 3655
rect 16850 3652 16856 3664
rect 16347 3624 16856 3652
rect 16347 3621 16359 3624
rect 16301 3615 16359 3621
rect 16850 3612 16856 3624
rect 16908 3612 16914 3664
rect 17589 3655 17647 3661
rect 17589 3621 17601 3655
rect 17635 3652 17647 3655
rect 19150 3652 19156 3664
rect 17635 3624 19156 3652
rect 17635 3621 17647 3624
rect 17589 3615 17647 3621
rect 19150 3612 19156 3624
rect 19208 3612 19214 3664
rect 19334 3612 19340 3664
rect 19392 3652 19398 3664
rect 19429 3655 19487 3661
rect 19429 3652 19441 3655
rect 19392 3624 19441 3652
rect 19392 3612 19398 3624
rect 19429 3621 19441 3624
rect 19475 3621 19487 3655
rect 19429 3615 19487 3621
rect 31018 3612 31024 3664
rect 31076 3652 31082 3664
rect 31665 3655 31723 3661
rect 31665 3652 31677 3655
rect 31076 3624 31677 3652
rect 31076 3612 31082 3624
rect 31665 3621 31677 3624
rect 31711 3621 31723 3655
rect 31665 3615 31723 3621
rect 16945 3587 17003 3593
rect 16945 3553 16957 3587
rect 16991 3584 17003 3587
rect 17770 3584 17776 3596
rect 16991 3556 17776 3584
rect 16991 3553 17003 3556
rect 16945 3547 17003 3553
rect 17770 3544 17776 3556
rect 17828 3544 17834 3596
rect 18877 3587 18935 3593
rect 18877 3553 18889 3587
rect 18923 3584 18935 3587
rect 22465 3587 22523 3593
rect 22465 3584 22477 3587
rect 18923 3556 22477 3584
rect 18923 3553 18935 3556
rect 18877 3547 18935 3553
rect 22465 3553 22477 3556
rect 22511 3553 22523 3587
rect 22738 3584 22744 3596
rect 22699 3556 22744 3584
rect 22465 3547 22523 3553
rect 22738 3544 22744 3556
rect 22796 3544 22802 3596
rect 28534 3584 28540 3596
rect 28495 3556 28540 3584
rect 28534 3544 28540 3556
rect 28592 3544 28598 3596
rect 28813 3587 28871 3593
rect 28813 3553 28825 3587
rect 28859 3584 28871 3587
rect 30190 3584 30196 3596
rect 28859 3556 30196 3584
rect 28859 3553 28871 3556
rect 28813 3547 28871 3553
rect 30190 3544 30196 3556
rect 30248 3544 30254 3596
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 4249 3519 4307 3525
rect 4249 3516 4261 3519
rect 4212 3488 4261 3516
rect 4212 3476 4218 3488
rect 4249 3485 4261 3488
rect 4295 3485 4307 3519
rect 5166 3516 5172 3528
rect 5127 3488 5172 3516
rect 4249 3479 4307 3485
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 5994 3516 6000 3528
rect 5955 3488 6000 3516
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 6822 3516 6828 3528
rect 6783 3488 6828 3516
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 7650 3516 7656 3528
rect 7611 3488 7656 3516
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 8478 3516 8484 3528
rect 8439 3488 8484 3516
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 9306 3516 9312 3528
rect 9267 3488 9312 3516
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 10134 3516 10140 3528
rect 10095 3488 10140 3516
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 10962 3516 10968 3528
rect 10923 3488 10968 3516
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11701 3519 11759 3525
rect 11701 3485 11713 3519
rect 11747 3516 11759 3519
rect 11790 3516 11796 3528
rect 11747 3488 11796 3516
rect 11747 3485 11759 3488
rect 11701 3479 11759 3485
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 12345 3519 12403 3525
rect 12345 3485 12357 3519
rect 12391 3516 12403 3519
rect 12526 3516 12532 3528
rect 12391 3488 12532 3516
rect 12391 3485 12403 3488
rect 12345 3479 12403 3485
rect 12526 3476 12532 3488
rect 12584 3476 12590 3528
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3516 13047 3519
rect 13078 3516 13084 3528
rect 13035 3488 13084 3516
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 13630 3516 13636 3528
rect 13591 3488 13636 3516
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 15010 3516 15016 3528
rect 14971 3488 15016 3516
rect 15010 3476 15016 3488
rect 15068 3476 15074 3528
rect 15657 3519 15715 3525
rect 15657 3485 15669 3519
rect 15703 3516 15715 3519
rect 16390 3516 16396 3528
rect 15703 3488 16396 3516
rect 15703 3485 15715 3488
rect 15657 3479 15715 3485
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 21542 3516 21548 3528
rect 21503 3488 21548 3516
rect 21542 3476 21548 3488
rect 21600 3476 21606 3528
rect 25409 3519 25467 3525
rect 25409 3485 25421 3519
rect 25455 3516 25467 3519
rect 25498 3516 25504 3528
rect 25455 3488 25504 3516
rect 25455 3485 25467 3488
rect 25409 3479 25467 3485
rect 25498 3476 25504 3488
rect 25556 3476 25562 3528
rect 26510 3516 26516 3528
rect 26471 3488 26516 3516
rect 26510 3476 26516 3488
rect 26568 3476 26574 3528
rect 29730 3516 29736 3528
rect 29691 3488 29736 3516
rect 29730 3476 29736 3488
rect 29788 3476 29794 3528
rect 29914 3476 29920 3528
rect 29972 3516 29978 3528
rect 30377 3519 30435 3525
rect 30377 3516 30389 3519
rect 29972 3488 30389 3516
rect 29972 3476 29978 3488
rect 30377 3485 30389 3488
rect 30423 3485 30435 3519
rect 30377 3479 30435 3485
rect 30466 3476 30472 3528
rect 30524 3516 30530 3528
rect 31021 3519 31079 3525
rect 31021 3516 31033 3519
rect 30524 3488 31033 3516
rect 30524 3476 30530 3488
rect 31021 3485 31033 3488
rect 31067 3485 31079 3519
rect 31021 3479 31079 3485
rect 31846 3476 31852 3528
rect 31904 3516 31910 3528
rect 32309 3519 32367 3525
rect 32309 3516 32321 3519
rect 31904 3488 32321 3516
rect 31904 3476 31910 3488
rect 32309 3485 32321 3488
rect 32355 3485 32367 3519
rect 32309 3479 32367 3485
rect 32674 3476 32680 3528
rect 32732 3516 32738 3528
rect 32953 3519 33011 3525
rect 32953 3516 32965 3519
rect 32732 3488 32965 3516
rect 32732 3476 32738 3488
rect 32953 3485 32965 3488
rect 32999 3485 33011 3519
rect 32953 3479 33011 3485
rect 33226 3476 33232 3528
rect 33284 3516 33290 3528
rect 33597 3519 33655 3525
rect 33597 3516 33609 3519
rect 33284 3488 33609 3516
rect 33284 3476 33290 3488
rect 33597 3485 33609 3488
rect 33643 3485 33655 3519
rect 33597 3479 33655 3485
rect 35161 3519 35219 3525
rect 35161 3485 35173 3519
rect 35207 3516 35219 3519
rect 35342 3516 35348 3528
rect 35207 3488 35348 3516
rect 35207 3485 35219 3488
rect 35161 3479 35219 3485
rect 35342 3476 35348 3488
rect 35400 3476 35406 3528
rect 35434 3476 35440 3528
rect 35492 3516 35498 3528
rect 35621 3519 35679 3525
rect 35621 3516 35633 3519
rect 35492 3488 35633 3516
rect 35492 3476 35498 3488
rect 35621 3485 35633 3488
rect 35667 3485 35679 3519
rect 36262 3516 36268 3528
rect 36223 3488 36268 3516
rect 35621 3479 35679 3485
rect 36262 3476 36268 3488
rect 36320 3476 36326 3528
rect 37090 3516 37096 3528
rect 37051 3488 37096 3516
rect 37090 3476 37096 3488
rect 37148 3476 37154 3528
rect 37918 3516 37924 3528
rect 37879 3488 37924 3516
rect 37918 3476 37924 3488
rect 37976 3476 37982 3528
rect 39022 3516 39028 3528
rect 38983 3488 39028 3516
rect 39022 3476 39028 3488
rect 39080 3476 39086 3528
rect 40402 3516 40408 3528
rect 40363 3488 40408 3516
rect 40402 3476 40408 3488
rect 40460 3476 40466 3528
rect 40865 3519 40923 3525
rect 40865 3485 40877 3519
rect 40911 3516 40923 3519
rect 40954 3516 40960 3528
rect 40911 3488 40960 3516
rect 40911 3485 40923 3488
rect 40865 3479 40923 3485
rect 40954 3476 40960 3488
rect 41012 3476 41018 3528
rect 41506 3516 41512 3528
rect 41467 3488 41512 3516
rect 41506 3476 41512 3488
rect 41564 3476 41570 3528
rect 42886 3516 42892 3528
rect 42847 3488 42892 3516
rect 42886 3476 42892 3488
rect 42944 3476 42950 3528
rect 43162 3476 43168 3528
rect 43220 3516 43226 3528
rect 43349 3519 43407 3525
rect 43349 3516 43361 3519
rect 43220 3488 43361 3516
rect 43220 3476 43226 3488
rect 43349 3485 43361 3488
rect 43395 3485 43407 3519
rect 43349 3479 43407 3485
rect 44818 3476 44824 3528
rect 44876 3516 44882 3528
rect 45189 3519 45247 3525
rect 45189 3516 45201 3519
rect 44876 3488 45201 3516
rect 44876 3476 44882 3488
rect 45189 3485 45201 3488
rect 45235 3485 45247 3519
rect 45189 3479 45247 3485
rect 45646 3476 45652 3528
rect 45704 3516 45710 3528
rect 45833 3519 45891 3525
rect 45833 3516 45845 3519
rect 45704 3488 45845 3516
rect 45704 3476 45710 3488
rect 45833 3485 45845 3488
rect 45879 3485 45891 3519
rect 46474 3516 46480 3528
rect 46435 3488 46480 3516
rect 45833 3479 45891 3485
rect 46474 3476 46480 3488
rect 46532 3476 46538 3528
rect 46750 3476 46756 3528
rect 46808 3516 46814 3528
rect 47121 3519 47179 3525
rect 47121 3516 47133 3519
rect 46808 3488 47133 3516
rect 46808 3476 46814 3488
rect 47121 3485 47133 3488
rect 47167 3485 47179 3519
rect 47121 3479 47179 3485
rect 47302 3476 47308 3528
rect 47360 3516 47366 3528
rect 47765 3519 47823 3525
rect 47765 3516 47777 3519
rect 47360 3488 47777 3516
rect 47360 3476 47366 3488
rect 47765 3485 47777 3488
rect 47811 3485 47823 3519
rect 47765 3479 47823 3485
rect 18874 3408 18880 3460
rect 18932 3448 18938 3460
rect 20073 3451 20131 3457
rect 20073 3448 20085 3451
rect 18932 3420 20085 3448
rect 18932 3408 18938 3420
rect 20073 3417 20085 3420
rect 20119 3417 20131 3451
rect 20073 3411 20131 3417
rect 20162 3408 20168 3460
rect 20220 3448 20226 3460
rect 21085 3451 21143 3457
rect 20220 3420 20265 3448
rect 20220 3408 20226 3420
rect 21085 3417 21097 3451
rect 21131 3448 21143 3451
rect 21358 3448 21364 3460
rect 21131 3420 21364 3448
rect 21131 3417 21143 3420
rect 21085 3411 21143 3417
rect 21358 3408 21364 3420
rect 21416 3408 21422 3460
rect 22557 3451 22615 3457
rect 22557 3417 22569 3451
rect 22603 3417 22615 3451
rect 28718 3448 28724 3460
rect 28679 3420 28724 3448
rect 22557 3411 22615 3417
rect 21821 3383 21879 3389
rect 21821 3349 21833 3383
rect 21867 3380 21879 3383
rect 22572 3380 22600 3411
rect 28718 3408 28724 3420
rect 28776 3408 28782 3460
rect 29638 3408 29644 3460
rect 29696 3448 29702 3460
rect 30834 3448 30840 3460
rect 29696 3420 30840 3448
rect 29696 3408 29702 3420
rect 30834 3408 30840 3420
rect 30892 3408 30898 3460
rect 25406 3380 25412 3392
rect 21867 3352 22600 3380
rect 25367 3352 25412 3380
rect 21867 3349 21879 3352
rect 21821 3343 21879 3349
rect 25406 3340 25412 3352
rect 25464 3340 25470 3392
rect 26697 3383 26755 3389
rect 26697 3349 26709 3383
rect 26743 3380 26755 3383
rect 28074 3380 28080 3392
rect 26743 3352 28080 3380
rect 26743 3349 26755 3352
rect 26697 3343 26755 3349
rect 28074 3340 28080 3352
rect 28132 3340 28138 3392
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 20073 3179 20131 3185
rect 20073 3145 20085 3179
rect 20119 3176 20131 3179
rect 20162 3176 20168 3188
rect 20119 3148 20168 3176
rect 20119 3145 20131 3148
rect 20073 3139 20131 3145
rect 20162 3136 20168 3148
rect 20220 3136 20226 3188
rect 20530 3108 20536 3120
rect 18248 3080 20536 3108
rect 18248 3049 18276 3080
rect 20530 3068 20536 3080
rect 20588 3068 20594 3120
rect 22186 3108 22192 3120
rect 22147 3080 22192 3108
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 23750 3068 23756 3120
rect 23808 3108 23814 3120
rect 23845 3111 23903 3117
rect 23845 3108 23857 3111
rect 23808 3080 23857 3108
rect 23808 3068 23814 3080
rect 23845 3077 23857 3080
rect 23891 3077 23903 3111
rect 25406 3108 25412 3120
rect 25367 3080 25412 3108
rect 23845 3071 23903 3077
rect 25406 3068 25412 3080
rect 25464 3068 25470 3120
rect 28074 3108 28080 3120
rect 28035 3080 28080 3108
rect 28074 3068 28080 3080
rect 28132 3068 28138 3120
rect 29641 3111 29699 3117
rect 29641 3077 29653 3111
rect 29687 3108 29699 3111
rect 30285 3111 30343 3117
rect 30285 3108 30297 3111
rect 29687 3080 30297 3108
rect 29687 3077 29699 3080
rect 29641 3071 29699 3077
rect 30285 3077 30297 3080
rect 30331 3077 30343 3111
rect 30285 3071 30343 3077
rect 18233 3043 18291 3049
rect 18233 3009 18245 3043
rect 18279 3009 18291 3043
rect 18874 3040 18880 3052
rect 18835 3012 18880 3040
rect 18233 3003 18291 3009
rect 18874 3000 18880 3012
rect 18932 3000 18938 3052
rect 20346 3040 20352 3052
rect 20307 3012 20352 3040
rect 20346 3000 20352 3012
rect 20404 3000 20410 3052
rect 21361 3043 21419 3049
rect 21361 3009 21373 3043
rect 21407 3040 21419 3043
rect 21542 3040 21548 3052
rect 21407 3012 21548 3040
rect 21407 3009 21419 3012
rect 21361 3003 21419 3009
rect 21542 3000 21548 3012
rect 21600 3000 21606 3052
rect 30098 3000 30104 3052
rect 30156 3040 30162 3052
rect 30377 3043 30435 3049
rect 30377 3040 30389 3043
rect 30156 3012 30389 3040
rect 30156 3000 30162 3012
rect 30377 3009 30389 3012
rect 30423 3009 30435 3043
rect 30377 3003 30435 3009
rect 4709 2975 4767 2981
rect 4709 2941 4721 2975
rect 4755 2972 4767 2975
rect 5442 2972 5448 2984
rect 4755 2944 5448 2972
rect 4755 2941 4767 2944
rect 4709 2935 4767 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 7285 2975 7343 2981
rect 7285 2941 7297 2975
rect 7331 2972 7343 2975
rect 7926 2972 7932 2984
rect 7331 2944 7932 2972
rect 7331 2941 7343 2944
rect 7285 2935 7343 2941
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2972 9275 2975
rect 9858 2972 9864 2984
rect 9263 2944 9864 2972
rect 9263 2941 9275 2944
rect 9217 2935 9275 2941
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 14369 2975 14427 2981
rect 14369 2941 14381 2975
rect 14415 2972 14427 2975
rect 15286 2972 15292 2984
rect 14415 2944 15292 2972
rect 14415 2941 14427 2944
rect 14369 2935 14427 2941
rect 15286 2932 15292 2944
rect 15344 2932 15350 2984
rect 15657 2975 15715 2981
rect 15657 2941 15669 2975
rect 15703 2972 15715 2975
rect 17494 2972 17500 2984
rect 15703 2944 17500 2972
rect 15703 2941 15715 2944
rect 15657 2935 15715 2941
rect 17494 2932 17500 2944
rect 17552 2932 17558 2984
rect 17589 2975 17647 2981
rect 17589 2941 17601 2975
rect 17635 2972 17647 2975
rect 17635 2944 19288 2972
rect 17635 2941 17647 2944
rect 17589 2935 17647 2941
rect 4065 2907 4123 2913
rect 4065 2873 4077 2907
rect 4111 2904 4123 2907
rect 4890 2904 4896 2916
rect 4111 2876 4896 2904
rect 4111 2873 4123 2876
rect 4065 2867 4123 2873
rect 4890 2864 4896 2876
rect 4948 2864 4954 2916
rect 5353 2907 5411 2913
rect 5353 2873 5365 2907
rect 5399 2904 5411 2907
rect 6270 2904 6276 2916
rect 5399 2876 6276 2904
rect 5399 2873 5411 2876
rect 5353 2867 5411 2873
rect 6270 2864 6276 2876
rect 6328 2864 6334 2916
rect 8754 2904 8760 2916
rect 7944 2876 8760 2904
rect 2777 2839 2835 2845
rect 2777 2805 2789 2839
rect 2823 2836 2835 2839
rect 3142 2836 3148 2848
rect 2823 2808 3148 2836
rect 2823 2805 2835 2808
rect 2777 2799 2835 2805
rect 3142 2796 3148 2808
rect 3200 2796 3206 2848
rect 3421 2839 3479 2845
rect 3421 2805 3433 2839
rect 3467 2836 3479 2839
rect 3878 2836 3884 2848
rect 3467 2808 3884 2836
rect 3467 2805 3479 2808
rect 3421 2799 3479 2805
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 5997 2839 6055 2845
rect 5997 2805 6009 2839
rect 6043 2836 6055 2839
rect 6546 2836 6552 2848
rect 6043 2808 6552 2836
rect 6043 2805 6055 2808
rect 5997 2799 6055 2805
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 7944 2845 7972 2876
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 10505 2907 10563 2913
rect 10505 2873 10517 2907
rect 10551 2904 10563 2907
rect 11238 2904 11244 2916
rect 10551 2876 11244 2904
rect 10551 2873 10563 2876
rect 10505 2867 10563 2873
rect 11238 2864 11244 2876
rect 11296 2864 11302 2916
rect 12437 2907 12495 2913
rect 12437 2873 12449 2907
rect 12483 2904 12495 2907
rect 13354 2904 13360 2916
rect 12483 2876 13360 2904
rect 12483 2873 12495 2876
rect 12437 2867 12495 2873
rect 13354 2864 13360 2876
rect 13412 2864 13418 2916
rect 13725 2907 13783 2913
rect 13725 2873 13737 2907
rect 13771 2904 13783 2907
rect 14458 2904 14464 2916
rect 13771 2876 14464 2904
rect 13771 2873 13783 2876
rect 13725 2867 13783 2873
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 16301 2907 16359 2913
rect 16301 2873 16313 2907
rect 16347 2904 16359 2907
rect 18046 2904 18052 2916
rect 16347 2876 18052 2904
rect 16347 2873 16359 2876
rect 16301 2867 16359 2873
rect 18046 2864 18052 2876
rect 18104 2864 18110 2916
rect 7929 2839 7987 2845
rect 7929 2805 7941 2839
rect 7975 2805 7987 2839
rect 7929 2799 7987 2805
rect 8573 2839 8631 2845
rect 8573 2805 8585 2839
rect 8619 2836 8631 2839
rect 9030 2836 9036 2848
rect 8619 2808 9036 2836
rect 8619 2805 8631 2808
rect 8573 2799 8631 2805
rect 9030 2796 9036 2808
rect 9088 2796 9094 2848
rect 9861 2839 9919 2845
rect 9861 2805 9873 2839
rect 9907 2836 9919 2839
rect 10686 2836 10692 2848
rect 9907 2808 10692 2836
rect 9907 2805 9919 2808
rect 9861 2799 9919 2805
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 11149 2839 11207 2845
rect 11149 2805 11161 2839
rect 11195 2836 11207 2839
rect 12066 2836 12072 2848
rect 11195 2808 12072 2836
rect 11195 2805 11207 2808
rect 11149 2799 11207 2805
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 13081 2839 13139 2845
rect 13081 2805 13093 2839
rect 13127 2836 13139 2839
rect 13906 2836 13912 2848
rect 13127 2808 13912 2836
rect 13127 2805 13139 2808
rect 13081 2799 13139 2805
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 15013 2839 15071 2845
rect 15013 2805 15025 2839
rect 15059 2836 15071 2839
rect 15838 2836 15844 2848
rect 15059 2808 15844 2836
rect 15059 2805 15071 2808
rect 15013 2799 15071 2805
rect 15838 2796 15844 2808
rect 15896 2796 15902 2848
rect 19260 2836 19288 2944
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 22097 2975 22155 2981
rect 22097 2972 22109 2975
rect 19392 2944 22109 2972
rect 19392 2932 19398 2944
rect 22097 2941 22109 2944
rect 22143 2941 22155 2975
rect 22462 2972 22468 2984
rect 22423 2944 22468 2972
rect 22097 2935 22155 2941
rect 22462 2932 22468 2944
rect 22520 2932 22526 2984
rect 23753 2975 23811 2981
rect 23753 2941 23765 2975
rect 23799 2941 23811 2975
rect 24394 2972 24400 2984
rect 24355 2944 24400 2972
rect 23753 2935 23811 2941
rect 19521 2907 19579 2913
rect 19521 2873 19533 2907
rect 19567 2904 19579 2907
rect 23768 2904 23796 2935
rect 24394 2932 24400 2944
rect 24452 2932 24458 2984
rect 24578 2932 24584 2984
rect 24636 2972 24642 2984
rect 25317 2975 25375 2981
rect 25317 2972 25329 2975
rect 24636 2944 25329 2972
rect 24636 2932 24642 2944
rect 25317 2941 25329 2944
rect 25363 2941 25375 2975
rect 25774 2972 25780 2984
rect 25735 2944 25780 2972
rect 25317 2935 25375 2941
rect 25774 2932 25780 2944
rect 25832 2932 25838 2984
rect 27154 2972 27160 2984
rect 27115 2944 27160 2972
rect 27154 2932 27160 2944
rect 27212 2932 27218 2984
rect 28169 2975 28227 2981
rect 28169 2941 28181 2975
rect 28215 2972 28227 2975
rect 29178 2972 29184 2984
rect 28215 2944 29184 2972
rect 28215 2941 28227 2944
rect 28169 2935 28227 2941
rect 29178 2932 29184 2944
rect 29236 2932 29242 2984
rect 29362 2972 29368 2984
rect 29323 2944 29368 2972
rect 29362 2932 29368 2944
rect 29420 2932 29426 2984
rect 29733 2975 29791 2981
rect 29733 2941 29745 2975
rect 29779 2972 29791 2975
rect 31202 2972 31208 2984
rect 29779 2944 31208 2972
rect 29779 2941 29791 2944
rect 29733 2935 29791 2941
rect 31202 2932 31208 2944
rect 31260 2932 31266 2984
rect 32950 2932 32956 2984
rect 33008 2972 33014 2984
rect 33597 2975 33655 2981
rect 33597 2972 33609 2975
rect 33008 2944 33609 2972
rect 33008 2932 33014 2944
rect 33597 2941 33609 2944
rect 33643 2941 33655 2975
rect 33597 2935 33655 2941
rect 38746 2932 38752 2984
rect 38804 2972 38810 2984
rect 39393 2975 39451 2981
rect 39393 2972 39405 2975
rect 38804 2944 39405 2972
rect 38804 2932 38810 2944
rect 39393 2941 39405 2944
rect 39439 2941 39451 2975
rect 39393 2935 39451 2941
rect 40678 2932 40684 2984
rect 40736 2972 40742 2984
rect 41325 2975 41383 2981
rect 41325 2972 41337 2975
rect 40736 2944 41337 2972
rect 40736 2932 40742 2944
rect 41325 2941 41337 2944
rect 41371 2941 41383 2975
rect 41325 2935 41383 2941
rect 42610 2932 42616 2984
rect 42668 2972 42674 2984
rect 43257 2975 43315 2981
rect 43257 2972 43269 2975
rect 42668 2944 43269 2972
rect 42668 2932 42674 2944
rect 43257 2941 43269 2944
rect 43303 2941 43315 2975
rect 43257 2935 43315 2941
rect 44542 2932 44548 2984
rect 44600 2972 44606 2984
rect 45189 2975 45247 2981
rect 45189 2972 45201 2975
rect 44600 2944 45201 2972
rect 44600 2932 44606 2944
rect 45189 2941 45201 2944
rect 45235 2941 45247 2975
rect 45189 2935 45247 2941
rect 19567 2876 23796 2904
rect 19567 2873 19579 2876
rect 19521 2867 19579 2873
rect 34790 2864 34796 2916
rect 34848 2904 34854 2916
rect 35529 2907 35587 2913
rect 35529 2904 35541 2907
rect 34848 2876 35541 2904
rect 34848 2864 34854 2876
rect 35529 2873 35541 2876
rect 35575 2873 35587 2907
rect 35529 2867 35587 2873
rect 19978 2836 19984 2848
rect 19260 2808 19984 2836
rect 19978 2796 19984 2808
rect 20036 2796 20042 2848
rect 21361 2839 21419 2845
rect 21361 2805 21373 2839
rect 21407 2836 21419 2839
rect 22830 2836 22836 2848
rect 21407 2808 22836 2836
rect 21407 2805 21419 2808
rect 21361 2799 21419 2805
rect 22830 2796 22836 2808
rect 22888 2796 22894 2848
rect 30190 2796 30196 2848
rect 30248 2836 30254 2848
rect 31113 2839 31171 2845
rect 31113 2836 31125 2839
rect 30248 2808 31125 2836
rect 30248 2796 30254 2808
rect 31113 2805 31125 2808
rect 31159 2805 31171 2839
rect 31113 2799 31171 2805
rect 31294 2796 31300 2848
rect 31352 2836 31358 2848
rect 32309 2839 32367 2845
rect 32309 2836 32321 2839
rect 31352 2808 32321 2836
rect 31352 2796 31358 2808
rect 32309 2805 32321 2808
rect 32355 2805 32367 2839
rect 32309 2799 32367 2805
rect 32398 2796 32404 2848
rect 32456 2836 32462 2848
rect 32953 2839 33011 2845
rect 32953 2836 32965 2839
rect 32456 2808 32965 2836
rect 32456 2796 32462 2808
rect 32953 2805 32965 2808
rect 32999 2805 33011 2839
rect 32953 2799 33011 2805
rect 33778 2796 33784 2848
rect 33836 2836 33842 2848
rect 34241 2839 34299 2845
rect 34241 2836 34253 2839
rect 33836 2808 34253 2836
rect 33836 2796 33842 2808
rect 34241 2805 34253 2808
rect 34287 2805 34299 2839
rect 34241 2799 34299 2805
rect 34330 2796 34336 2848
rect 34388 2836 34394 2848
rect 34885 2839 34943 2845
rect 34885 2836 34897 2839
rect 34388 2808 34897 2836
rect 34388 2796 34394 2808
rect 34885 2805 34897 2808
rect 34931 2805 34943 2839
rect 34885 2799 34943 2805
rect 35710 2796 35716 2848
rect 35768 2836 35774 2848
rect 36173 2839 36231 2845
rect 36173 2836 36185 2839
rect 35768 2808 36185 2836
rect 35768 2796 35774 2808
rect 36173 2805 36185 2808
rect 36219 2805 36231 2839
rect 36173 2799 36231 2805
rect 36814 2796 36820 2848
rect 36872 2836 36878 2848
rect 37461 2839 37519 2845
rect 37461 2836 37473 2839
rect 36872 2808 37473 2836
rect 36872 2796 36878 2808
rect 37461 2805 37473 2808
rect 37507 2805 37519 2839
rect 37461 2799 37519 2805
rect 37642 2796 37648 2848
rect 37700 2836 37706 2848
rect 38105 2839 38163 2845
rect 38105 2836 38117 2839
rect 37700 2808 38117 2836
rect 37700 2796 37706 2808
rect 38105 2805 38117 2808
rect 38151 2805 38163 2839
rect 38105 2799 38163 2805
rect 38194 2796 38200 2848
rect 38252 2836 38258 2848
rect 38749 2839 38807 2845
rect 38749 2836 38761 2839
rect 38252 2808 38761 2836
rect 38252 2796 38258 2808
rect 38749 2805 38761 2808
rect 38795 2805 38807 2839
rect 38749 2799 38807 2805
rect 39574 2796 39580 2848
rect 39632 2836 39638 2848
rect 40037 2839 40095 2845
rect 40037 2836 40049 2839
rect 39632 2808 40049 2836
rect 39632 2796 39638 2808
rect 40037 2805 40049 2808
rect 40083 2805 40095 2839
rect 40037 2799 40095 2805
rect 40126 2796 40132 2848
rect 40184 2836 40190 2848
rect 40681 2839 40739 2845
rect 40681 2836 40693 2839
rect 40184 2808 40693 2836
rect 40184 2796 40190 2808
rect 40681 2805 40693 2808
rect 40727 2805 40739 2839
rect 40681 2799 40739 2805
rect 42058 2796 42064 2848
rect 42116 2836 42122 2848
rect 42613 2839 42671 2845
rect 42613 2836 42625 2839
rect 42116 2808 42625 2836
rect 42116 2796 42122 2808
rect 42613 2805 42625 2808
rect 42659 2805 42671 2839
rect 42613 2799 42671 2805
rect 43438 2796 43444 2848
rect 43496 2836 43502 2848
rect 43901 2839 43959 2845
rect 43901 2836 43913 2839
rect 43496 2808 43913 2836
rect 43496 2796 43502 2808
rect 43901 2805 43913 2808
rect 43947 2805 43959 2839
rect 43901 2799 43959 2805
rect 43990 2796 43996 2848
rect 44048 2836 44054 2848
rect 44545 2839 44603 2845
rect 44545 2836 44557 2839
rect 44048 2808 44557 2836
rect 44048 2796 44054 2808
rect 44545 2805 44557 2808
rect 44591 2805 44603 2839
rect 44545 2799 44603 2805
rect 45370 2796 45376 2848
rect 45428 2836 45434 2848
rect 45833 2839 45891 2845
rect 45833 2836 45845 2839
rect 45428 2808 45845 2836
rect 45428 2796 45434 2808
rect 45833 2805 45845 2808
rect 45879 2805 45891 2839
rect 45833 2799 45891 2805
rect 45922 2796 45928 2848
rect 45980 2836 45986 2848
rect 46477 2839 46535 2845
rect 46477 2836 46489 2839
rect 45980 2808 46489 2836
rect 45980 2796 45986 2808
rect 46477 2805 46489 2808
rect 46523 2805 46535 2839
rect 46477 2799 46535 2805
rect 47026 2796 47032 2848
rect 47084 2836 47090 2848
rect 47765 2839 47823 2845
rect 47765 2836 47777 2839
rect 47084 2808 47777 2836
rect 47084 2796 47090 2808
rect 47765 2805 47777 2808
rect 47811 2805 47823 2839
rect 47765 2799 47823 2805
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 18877 2635 18935 2641
rect 18877 2601 18889 2635
rect 18923 2632 18935 2635
rect 19334 2632 19340 2644
rect 18923 2604 19340 2632
rect 18923 2601 18935 2604
rect 18877 2595 18935 2601
rect 19334 2592 19340 2604
rect 19392 2592 19398 2644
rect 21361 2635 21419 2641
rect 21361 2601 21373 2635
rect 21407 2632 21419 2635
rect 22186 2632 22192 2644
rect 21407 2604 22192 2632
rect 21407 2601 21419 2604
rect 21361 2595 21419 2601
rect 22186 2592 22192 2604
rect 22244 2592 22250 2644
rect 26418 2632 26424 2644
rect 26379 2604 26424 2632
rect 26418 2592 26424 2604
rect 26476 2592 26482 2644
rect 29178 2592 29184 2644
rect 29236 2632 29242 2644
rect 30561 2635 30619 2641
rect 30561 2632 30573 2635
rect 29236 2604 30573 2632
rect 29236 2592 29242 2604
rect 30561 2601 30573 2604
rect 30607 2601 30619 2635
rect 31202 2632 31208 2644
rect 31163 2604 31208 2632
rect 30561 2595 30619 2601
rect 31202 2592 31208 2604
rect 31260 2592 31266 2644
rect 5353 2567 5411 2573
rect 5353 2533 5365 2567
rect 5399 2564 5411 2567
rect 7098 2564 7104 2576
rect 5399 2536 7104 2564
rect 5399 2533 5411 2536
rect 5353 2527 5411 2533
rect 7098 2524 7104 2536
rect 7156 2524 7162 2576
rect 7929 2567 7987 2573
rect 7929 2533 7941 2567
rect 7975 2564 7987 2567
rect 9582 2564 9588 2576
rect 7975 2536 9588 2564
rect 7975 2533 7987 2536
rect 7929 2527 7987 2533
rect 9582 2524 9588 2536
rect 9640 2524 9646 2576
rect 9861 2567 9919 2573
rect 9861 2533 9873 2567
rect 9907 2564 9919 2567
rect 11514 2564 11520 2576
rect 9907 2536 11520 2564
rect 9907 2533 9919 2536
rect 9861 2527 9919 2533
rect 11514 2524 11520 2536
rect 11572 2524 11578 2576
rect 12437 2567 12495 2573
rect 12437 2533 12449 2567
rect 12483 2564 12495 2567
rect 14182 2564 14188 2576
rect 12483 2536 14188 2564
rect 12483 2533 12495 2536
rect 12437 2527 12495 2533
rect 14182 2524 14188 2536
rect 14240 2524 14246 2576
rect 17589 2567 17647 2573
rect 17589 2533 17601 2567
rect 17635 2564 17647 2567
rect 20254 2564 20260 2576
rect 17635 2536 20260 2564
rect 17635 2533 17647 2536
rect 17589 2527 17647 2533
rect 20254 2524 20260 2536
rect 20312 2524 20318 2576
rect 20625 2567 20683 2573
rect 20625 2533 20637 2567
rect 20671 2564 20683 2567
rect 20671 2536 24992 2564
rect 20671 2533 20683 2536
rect 20625 2527 20683 2533
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2496 2835 2499
rect 3510 2496 3516 2508
rect 2823 2468 3516 2496
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 3510 2456 3516 2468
rect 3568 2456 3574 2508
rect 7285 2499 7343 2505
rect 7285 2465 7297 2499
rect 7331 2496 7343 2499
rect 8202 2496 8208 2508
rect 7331 2468 8208 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2496 8631 2499
rect 10410 2496 10416 2508
rect 8619 2468 10416 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 10410 2456 10416 2468
rect 10468 2456 10474 2508
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2496 11207 2499
rect 12802 2496 12808 2508
rect 11195 2468 12808 2496
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 12802 2456 12808 2468
rect 12860 2456 12866 2508
rect 13081 2499 13139 2505
rect 13081 2465 13093 2499
rect 13127 2496 13139 2499
rect 14734 2496 14740 2508
rect 13127 2468 14740 2496
rect 13127 2465 13139 2468
rect 13081 2459 13139 2465
rect 14734 2456 14740 2468
rect 14792 2456 14798 2508
rect 15013 2499 15071 2505
rect 15013 2465 15025 2499
rect 15059 2496 15071 2499
rect 16666 2496 16672 2508
rect 15059 2468 16672 2496
rect 15059 2465 15071 2468
rect 15013 2459 15071 2465
rect 16666 2456 16672 2468
rect 16724 2456 16730 2508
rect 18874 2496 18880 2508
rect 17512 2468 18880 2496
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 2590 2428 2596 2440
rect 2179 2400 2596 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 4614 2428 4620 2440
rect 3467 2400 4620 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2428 4767 2431
rect 5718 2428 5724 2440
rect 4755 2400 5724 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 10505 2431 10563 2437
rect 6043 2400 6914 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6886 2360 6914 2400
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 12250 2428 12256 2440
rect 10551 2400 12256 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 12250 2388 12256 2400
rect 12308 2388 12314 2440
rect 13725 2431 13783 2437
rect 13725 2397 13737 2431
rect 13771 2428 13783 2431
rect 15562 2428 15568 2440
rect 13771 2400 15568 2428
rect 13771 2397 13783 2400
rect 13725 2391 13783 2397
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2397 15715 2431
rect 15657 2391 15715 2397
rect 16301 2431 16359 2437
rect 16301 2397 16313 2431
rect 16347 2428 16359 2431
rect 17512 2428 17540 2468
rect 18874 2456 18880 2468
rect 18932 2456 18938 2508
rect 19981 2499 20039 2505
rect 19981 2465 19993 2499
rect 20027 2496 20039 2499
rect 22741 2499 22799 2505
rect 22741 2496 22753 2499
rect 20027 2468 22753 2496
rect 20027 2465 20039 2468
rect 19981 2459 20039 2465
rect 22741 2465 22753 2468
rect 22787 2465 22799 2499
rect 23014 2496 23020 2508
rect 22975 2468 23020 2496
rect 22741 2459 22799 2465
rect 23014 2456 23020 2468
rect 23072 2456 23078 2508
rect 24964 2505 24992 2536
rect 32122 2524 32128 2576
rect 32180 2564 32186 2576
rect 33597 2567 33655 2573
rect 33597 2564 33609 2567
rect 32180 2536 33609 2564
rect 32180 2524 32186 2536
rect 33597 2533 33609 2536
rect 33643 2533 33655 2567
rect 33597 2527 33655 2533
rect 34606 2524 34612 2576
rect 34664 2564 34670 2576
rect 36173 2567 36231 2573
rect 36173 2564 36185 2567
rect 34664 2536 36185 2564
rect 34664 2524 34670 2536
rect 36173 2533 36185 2536
rect 36219 2533 36231 2567
rect 36173 2527 36231 2533
rect 38470 2524 38476 2576
rect 38528 2564 38534 2576
rect 40037 2567 40095 2573
rect 40037 2564 40049 2567
rect 38528 2536 40049 2564
rect 38528 2524 38534 2536
rect 40037 2533 40049 2536
rect 40083 2533 40095 2567
rect 40037 2527 40095 2533
rect 42334 2524 42340 2576
rect 42392 2564 42398 2576
rect 43901 2567 43959 2573
rect 43901 2564 43913 2567
rect 42392 2536 43913 2564
rect 42392 2524 42398 2536
rect 43901 2533 43913 2536
rect 43947 2533 43959 2567
rect 43901 2527 43959 2533
rect 45094 2524 45100 2576
rect 45152 2564 45158 2576
rect 46477 2567 46535 2573
rect 46477 2564 46489 2567
rect 45152 2536 46489 2564
rect 45152 2524 45158 2536
rect 46477 2533 46489 2536
rect 46523 2533 46535 2567
rect 46477 2527 46535 2533
rect 24949 2499 25007 2505
rect 24949 2465 24961 2499
rect 24995 2465 25007 2499
rect 25498 2496 25504 2508
rect 25459 2468 25504 2496
rect 24949 2459 25007 2465
rect 25498 2456 25504 2468
rect 25556 2456 25562 2508
rect 28258 2496 28264 2508
rect 28219 2468 28264 2496
rect 28258 2456 28264 2468
rect 28316 2456 28322 2508
rect 28629 2499 28687 2505
rect 28629 2465 28641 2499
rect 28675 2496 28687 2499
rect 29730 2496 29736 2508
rect 28675 2468 29736 2496
rect 28675 2465 28687 2468
rect 28629 2459 28687 2465
rect 29730 2456 29736 2468
rect 29788 2456 29794 2508
rect 31570 2456 31576 2508
rect 31628 2496 31634 2508
rect 32953 2499 33011 2505
rect 32953 2496 32965 2499
rect 31628 2468 32965 2496
rect 31628 2456 31634 2468
rect 32953 2465 32965 2468
rect 32999 2465 33011 2499
rect 32953 2459 33011 2465
rect 33502 2456 33508 2508
rect 33560 2496 33566 2508
rect 34885 2499 34943 2505
rect 34885 2496 34897 2499
rect 33560 2468 34897 2496
rect 33560 2456 33566 2468
rect 34885 2465 34897 2468
rect 34931 2465 34943 2499
rect 34885 2459 34943 2465
rect 36538 2456 36544 2508
rect 36596 2496 36602 2508
rect 38105 2499 38163 2505
rect 38105 2496 38117 2499
rect 36596 2468 38117 2496
rect 36596 2456 36602 2468
rect 38105 2465 38117 2468
rect 38151 2465 38163 2499
rect 38105 2459 38163 2465
rect 39298 2456 39304 2508
rect 39356 2496 39362 2508
rect 40681 2499 40739 2505
rect 40681 2496 40693 2499
rect 39356 2468 40693 2496
rect 39356 2456 39362 2468
rect 40681 2465 40693 2468
rect 40727 2465 40739 2499
rect 40681 2459 40739 2465
rect 41230 2456 41236 2508
rect 41288 2496 41294 2508
rect 42613 2499 42671 2505
rect 42613 2496 42625 2499
rect 41288 2468 42625 2496
rect 41288 2456 41294 2468
rect 42613 2465 42625 2468
rect 42659 2465 42671 2499
rect 42613 2459 42671 2465
rect 43714 2456 43720 2508
rect 43772 2496 43778 2508
rect 45189 2499 45247 2505
rect 45189 2496 45201 2499
rect 43772 2468 45201 2496
rect 43772 2456 43778 2468
rect 45189 2465 45201 2468
rect 45235 2465 45247 2499
rect 45189 2459 45247 2465
rect 16347 2400 17540 2428
rect 18233 2431 18291 2437
rect 16347 2397 16359 2400
rect 16301 2391 16359 2397
rect 18233 2397 18245 2431
rect 18279 2428 18291 2431
rect 20806 2428 20812 2440
rect 18279 2400 20812 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 7374 2360 7380 2372
rect 6886 2332 7380 2360
rect 7374 2320 7380 2332
rect 7432 2320 7438 2372
rect 15672 2360 15700 2391
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 21085 2431 21143 2437
rect 21085 2397 21097 2431
rect 21131 2397 21143 2431
rect 21085 2391 21143 2397
rect 22189 2431 22247 2437
rect 22189 2397 22201 2431
rect 22235 2428 22247 2431
rect 30098 2428 30104 2440
rect 22235 2400 22600 2428
rect 30059 2400 30104 2428
rect 22235 2397 22247 2400
rect 22189 2391 22247 2397
rect 18322 2360 18328 2372
rect 15672 2332 18328 2360
rect 18322 2320 18328 2332
rect 18380 2320 18386 2372
rect 20346 2320 20352 2372
rect 20404 2360 20410 2372
rect 21100 2360 21128 2391
rect 20404 2332 21128 2360
rect 20404 2320 20410 2332
rect 22572 2292 22600 2400
rect 30098 2388 30104 2400
rect 30156 2388 30162 2440
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 30800 2400 32321 2428
rect 30800 2388 30806 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 34054 2388 34060 2440
rect 34112 2428 34118 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 34112 2400 35541 2428
rect 34112 2388 34118 2400
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 35529 2391 35587 2397
rect 35986 2388 35992 2440
rect 36044 2428 36050 2440
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 36044 2400 37473 2428
rect 36044 2388 36050 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 38749 2431 38807 2437
rect 38749 2397 38761 2431
rect 38795 2397 38807 2431
rect 38749 2391 38807 2397
rect 22830 2320 22836 2372
rect 22888 2360 22894 2372
rect 25038 2360 25044 2372
rect 22888 2332 22933 2360
rect 24999 2332 25044 2360
rect 22888 2320 22894 2332
rect 25038 2320 25044 2332
rect 25096 2320 25102 2372
rect 28537 2363 28595 2369
rect 28537 2329 28549 2363
rect 28583 2329 28595 2363
rect 28537 2323 28595 2329
rect 24578 2292 24584 2304
rect 22572 2264 24584 2292
rect 24578 2252 24584 2264
rect 24636 2252 24642 2304
rect 28552 2292 28580 2323
rect 37366 2320 37372 2372
rect 37424 2360 37430 2372
rect 38764 2360 38792 2391
rect 39850 2388 39856 2440
rect 39908 2428 39914 2440
rect 41325 2431 41383 2437
rect 41325 2428 41337 2431
rect 39908 2400 41337 2428
rect 39908 2388 39914 2400
rect 41325 2397 41337 2400
rect 41371 2397 41383 2431
rect 41325 2391 41383 2397
rect 41782 2388 41788 2440
rect 41840 2428 41846 2440
rect 43257 2431 43315 2437
rect 43257 2428 43269 2431
rect 41840 2400 43269 2428
rect 41840 2388 41846 2400
rect 43257 2397 43269 2400
rect 43303 2397 43315 2431
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 43257 2391 43315 2397
rect 45526 2400 45845 2428
rect 37424 2332 38792 2360
rect 37424 2320 37430 2332
rect 44266 2320 44272 2372
rect 44324 2360 44330 2372
rect 45526 2360 45554 2400
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 46198 2388 46204 2440
rect 46256 2428 46262 2440
rect 47765 2431 47823 2437
rect 47765 2428 47777 2431
rect 46256 2400 47777 2428
rect 46256 2388 46262 2400
rect 47765 2397 47777 2400
rect 47811 2397 47823 2431
rect 47765 2391 47823 2397
rect 44324 2332 45554 2360
rect 44324 2320 44330 2332
rect 29825 2295 29883 2301
rect 29825 2292 29837 2295
rect 28552 2264 29837 2292
rect 29825 2261 29837 2264
rect 29871 2261 29883 2295
rect 29825 2255 29883 2261
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
<< via1 >>
rect 19708 47744 19760 47796
rect 22376 47744 22428 47796
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 4712 47243 4764 47252
rect 4712 47209 4721 47243
rect 4721 47209 4755 47243
rect 4755 47209 4764 47243
rect 4712 47200 4764 47209
rect 5816 47200 5868 47252
rect 6000 47243 6052 47252
rect 6000 47209 6009 47243
rect 6009 47209 6043 47243
rect 6043 47209 6052 47243
rect 6000 47200 6052 47209
rect 7104 47243 7156 47252
rect 7104 47209 7113 47243
rect 7113 47209 7147 47243
rect 7147 47209 7156 47243
rect 7104 47200 7156 47209
rect 7748 47243 7800 47252
rect 7748 47209 7757 47243
rect 7757 47209 7791 47243
rect 7791 47209 7800 47243
rect 7748 47200 7800 47209
rect 8392 47243 8444 47252
rect 8392 47209 8401 47243
rect 8401 47209 8435 47243
rect 8435 47209 8444 47243
rect 8392 47200 8444 47209
rect 9128 47243 9180 47252
rect 9128 47209 9137 47243
rect 9137 47209 9171 47243
rect 9171 47209 9180 47243
rect 9128 47200 9180 47209
rect 10232 47243 10284 47252
rect 10232 47209 10241 47243
rect 10241 47209 10275 47243
rect 10275 47209 10284 47243
rect 10232 47200 10284 47209
rect 11152 47243 11204 47252
rect 11152 47209 11161 47243
rect 11161 47209 11195 47243
rect 11195 47209 11204 47243
rect 11152 47200 11204 47209
rect 12440 47243 12492 47252
rect 12440 47209 12449 47243
rect 12449 47209 12483 47243
rect 12483 47209 12492 47243
rect 13544 47243 13596 47252
rect 12440 47200 12492 47209
rect 13544 47209 13553 47243
rect 13553 47209 13587 47243
rect 13587 47209 13596 47243
rect 13544 47200 13596 47209
rect 16856 47200 16908 47252
rect 20168 47200 20220 47252
rect 20628 47243 20680 47252
rect 20628 47209 20637 47243
rect 20637 47209 20671 47243
rect 20671 47209 20680 47243
rect 20628 47200 20680 47209
rect 25688 47200 25740 47252
rect 26056 47243 26108 47252
rect 26056 47209 26065 47243
rect 26065 47209 26099 47243
rect 26099 47209 26108 47243
rect 26056 47200 26108 47209
rect 40408 47200 40460 47252
rect 44180 47200 44232 47252
rect 45928 47200 45980 47252
rect 19708 47132 19760 47184
rect 19892 47132 19944 47184
rect 10600 46860 10652 46912
rect 17132 46860 17184 46912
rect 18144 46928 18196 46980
rect 18696 46996 18748 47048
rect 19892 47039 19944 47048
rect 18972 46928 19024 46980
rect 19892 47005 19901 47039
rect 19901 47005 19935 47039
rect 19935 47005 19944 47039
rect 19892 46996 19944 47005
rect 20444 47039 20496 47048
rect 20444 47005 20453 47039
rect 20453 47005 20487 47039
rect 20487 47005 20496 47039
rect 20444 46996 20496 47005
rect 22100 47039 22152 47048
rect 22100 47005 22109 47039
rect 22109 47005 22143 47039
rect 22143 47005 22152 47039
rect 22100 46996 22152 47005
rect 25136 47039 25188 47048
rect 25136 47005 25145 47039
rect 25145 47005 25179 47039
rect 25179 47005 25188 47039
rect 25136 46996 25188 47005
rect 27804 47064 27856 47116
rect 25596 47039 25648 47048
rect 25596 47005 25605 47039
rect 25605 47005 25639 47039
rect 25639 47005 25648 47039
rect 25596 46996 25648 47005
rect 27712 47039 27764 47048
rect 27712 47005 27721 47039
rect 27721 47005 27755 47039
rect 27755 47005 27764 47039
rect 27712 46996 27764 47005
rect 30288 47064 30340 47116
rect 31208 47107 31260 47116
rect 31208 47073 31217 47107
rect 31217 47073 31251 47107
rect 31251 47073 31260 47107
rect 31208 47064 31260 47073
rect 33876 47132 33928 47184
rect 36360 47132 36412 47184
rect 36820 47132 36872 47184
rect 28908 47039 28960 47048
rect 26884 46928 26936 46980
rect 27160 46971 27212 46980
rect 27160 46937 27169 46971
rect 27169 46937 27203 46971
rect 27203 46937 27212 46971
rect 27160 46928 27212 46937
rect 18420 46860 18472 46912
rect 18604 46860 18656 46912
rect 21180 46860 21232 46912
rect 21456 46860 21508 46912
rect 24216 46860 24268 46912
rect 26424 46860 26476 46912
rect 28908 47005 28917 47039
rect 28917 47005 28951 47039
rect 28951 47005 28960 47039
rect 28908 46996 28960 47005
rect 30012 46996 30064 47048
rect 30840 46996 30892 47048
rect 31300 46996 31352 47048
rect 33692 47039 33744 47048
rect 30380 46928 30432 46980
rect 32036 46928 32088 46980
rect 33140 46928 33192 46980
rect 33692 47005 33701 47039
rect 33701 47005 33735 47039
rect 33735 47005 33744 47039
rect 33692 46996 33744 47005
rect 35532 47039 35584 47048
rect 29368 46860 29420 46912
rect 29828 46860 29880 46912
rect 34428 46928 34480 46980
rect 35532 47005 35541 47039
rect 35541 47005 35575 47039
rect 35575 47005 35584 47039
rect 35532 46996 35584 47005
rect 37648 47064 37700 47116
rect 38476 47132 38528 47184
rect 41788 47132 41840 47184
rect 44272 47132 44324 47184
rect 36360 47039 36412 47048
rect 36360 47005 36369 47039
rect 36369 47005 36403 47039
rect 36403 47005 36412 47039
rect 36360 46996 36412 47005
rect 37464 47039 37516 47048
rect 37464 47005 37473 47039
rect 37473 47005 37507 47039
rect 37507 47005 37516 47039
rect 37464 46996 37516 47005
rect 38384 47039 38436 47048
rect 38384 47005 38393 47039
rect 38393 47005 38427 47039
rect 38427 47005 38436 47039
rect 38384 46996 38436 47005
rect 38660 46996 38712 47048
rect 40224 46996 40276 47048
rect 36636 46928 36688 46980
rect 35532 46860 35584 46912
rect 35716 46860 35768 46912
rect 35992 46860 36044 46912
rect 37096 46860 37148 46912
rect 39396 46928 39448 46980
rect 37832 46860 37884 46912
rect 39948 46860 40000 46912
rect 40592 46903 40644 46912
rect 40592 46869 40601 46903
rect 40601 46869 40635 46903
rect 40635 46869 40644 46903
rect 40592 46860 40644 46869
rect 42432 46996 42484 47048
rect 43260 47039 43312 47048
rect 43260 47005 43269 47039
rect 43269 47005 43303 47039
rect 43303 47005 43312 47039
rect 43260 46996 43312 47005
rect 43904 46860 43956 46912
rect 44732 46860 44784 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 16120 46699 16172 46708
rect 16120 46665 16129 46699
rect 16129 46665 16163 46699
rect 16163 46665 16172 46699
rect 16120 46656 16172 46665
rect 17224 46656 17276 46708
rect 9496 46588 9548 46640
rect 6920 46563 6972 46572
rect 6920 46529 6929 46563
rect 6929 46529 6963 46563
rect 6963 46529 6972 46563
rect 6920 46520 6972 46529
rect 14648 46563 14700 46572
rect 14648 46529 14657 46563
rect 14657 46529 14691 46563
rect 14691 46529 14700 46563
rect 14648 46520 14700 46529
rect 15568 46563 15620 46572
rect 15568 46529 15577 46563
rect 15577 46529 15611 46563
rect 15611 46529 15620 46563
rect 15568 46520 15620 46529
rect 17408 46520 17460 46572
rect 18052 46520 18104 46572
rect 18328 46520 18380 46572
rect 18420 46563 18472 46572
rect 18420 46529 18429 46563
rect 18429 46529 18463 46563
rect 18463 46529 18472 46563
rect 21640 46656 21692 46708
rect 18972 46563 19024 46572
rect 18420 46520 18472 46529
rect 18972 46529 18981 46563
rect 18981 46529 19015 46563
rect 19015 46529 19024 46563
rect 18972 46520 19024 46529
rect 19984 46588 20036 46640
rect 19892 46520 19944 46572
rect 20444 46520 20496 46572
rect 21732 46588 21784 46640
rect 22100 46563 22152 46572
rect 22100 46529 22109 46563
rect 22109 46529 22143 46563
rect 22143 46529 22152 46563
rect 22836 46563 22888 46572
rect 22100 46520 22152 46529
rect 22836 46529 22845 46563
rect 22845 46529 22879 46563
rect 22879 46529 22888 46563
rect 22836 46520 22888 46529
rect 23848 46588 23900 46640
rect 30380 46656 30432 46708
rect 32680 46656 32732 46708
rect 34152 46656 34204 46708
rect 27160 46588 27212 46640
rect 27804 46631 27856 46640
rect 27804 46597 27813 46631
rect 27813 46597 27847 46631
rect 27847 46597 27856 46631
rect 27804 46588 27856 46597
rect 13912 46452 13964 46504
rect 17592 46452 17644 46504
rect 18604 46452 18656 46504
rect 19432 46452 19484 46504
rect 20904 46495 20956 46504
rect 20904 46461 20913 46495
rect 20913 46461 20947 46495
rect 20947 46461 20956 46495
rect 20904 46452 20956 46461
rect 21456 46495 21508 46504
rect 21456 46461 21469 46495
rect 21469 46461 21503 46495
rect 21503 46461 21508 46495
rect 24124 46563 24176 46572
rect 24124 46529 24133 46563
rect 24133 46529 24167 46563
rect 24167 46529 24176 46563
rect 24308 46563 24360 46572
rect 24124 46520 24176 46529
rect 24308 46529 24317 46563
rect 24317 46529 24351 46563
rect 24351 46529 24360 46563
rect 24308 46520 24360 46529
rect 25596 46520 25648 46572
rect 26976 46520 27028 46572
rect 27068 46520 27120 46572
rect 31576 46588 31628 46640
rect 33508 46588 33560 46640
rect 33600 46588 33652 46640
rect 29092 46563 29144 46572
rect 29092 46529 29101 46563
rect 29101 46529 29135 46563
rect 29135 46529 29144 46563
rect 29092 46520 29144 46529
rect 29644 46563 29696 46572
rect 29644 46529 29653 46563
rect 29653 46529 29687 46563
rect 29687 46529 29696 46563
rect 29644 46520 29696 46529
rect 30472 46563 30524 46572
rect 30472 46529 30481 46563
rect 30481 46529 30515 46563
rect 30515 46529 30524 46563
rect 30472 46520 30524 46529
rect 31300 46563 31352 46572
rect 31300 46529 31309 46563
rect 31309 46529 31343 46563
rect 31343 46529 31352 46563
rect 31300 46520 31352 46529
rect 33140 46520 33192 46572
rect 33232 46563 33284 46572
rect 33232 46529 33241 46563
rect 33241 46529 33275 46563
rect 33275 46529 33284 46563
rect 33232 46520 33284 46529
rect 26424 46495 26476 46504
rect 21456 46452 21508 46461
rect 15016 46384 15068 46436
rect 19340 46384 19392 46436
rect 22744 46384 22796 46436
rect 25412 46427 25464 46436
rect 25412 46393 25421 46427
rect 25421 46393 25455 46427
rect 25455 46393 25464 46427
rect 25412 46384 25464 46393
rect 26424 46461 26433 46495
rect 26433 46461 26467 46495
rect 26467 46461 26476 46495
rect 26424 46452 26476 46461
rect 26792 46452 26844 46504
rect 30932 46452 30984 46504
rect 31116 46495 31168 46504
rect 31116 46461 31125 46495
rect 31125 46461 31159 46495
rect 31159 46461 31168 46495
rect 31116 46452 31168 46461
rect 32312 46384 32364 46436
rect 37464 46656 37516 46708
rect 38200 46656 38252 46708
rect 41420 46656 41472 46708
rect 34428 46563 34480 46572
rect 34428 46529 34437 46563
rect 34437 46529 34471 46563
rect 34471 46529 34480 46563
rect 34428 46520 34480 46529
rect 34612 46563 34664 46572
rect 34612 46529 34621 46563
rect 34621 46529 34655 46563
rect 34655 46529 34664 46563
rect 34612 46520 34664 46529
rect 35348 46520 35400 46572
rect 35532 46520 35584 46572
rect 34796 46495 34848 46504
rect 34796 46461 34805 46495
rect 34805 46461 34839 46495
rect 34839 46461 34848 46495
rect 34796 46452 34848 46461
rect 36360 46452 36412 46504
rect 18788 46316 18840 46368
rect 19432 46359 19484 46368
rect 19432 46325 19441 46359
rect 19441 46325 19475 46359
rect 19475 46325 19484 46359
rect 19432 46316 19484 46325
rect 19984 46316 20036 46368
rect 24860 46316 24912 46368
rect 26240 46316 26292 46368
rect 33048 46316 33100 46368
rect 36268 46384 36320 46436
rect 36820 46588 36872 46640
rect 38476 46563 38528 46572
rect 36636 46495 36688 46504
rect 36636 46461 36645 46495
rect 36645 46461 36679 46495
rect 36679 46461 36688 46495
rect 36636 46452 36688 46461
rect 36912 46452 36964 46504
rect 38108 46452 38160 46504
rect 38476 46529 38485 46563
rect 38485 46529 38519 46563
rect 38519 46529 38528 46563
rect 38476 46520 38528 46529
rect 39580 46563 39632 46572
rect 38384 46452 38436 46504
rect 39580 46529 39589 46563
rect 39589 46529 39623 46563
rect 39623 46529 39632 46563
rect 39580 46520 39632 46529
rect 40224 46563 40276 46572
rect 40224 46529 40233 46563
rect 40233 46529 40267 46563
rect 40267 46529 40276 46563
rect 40224 46520 40276 46529
rect 40316 46520 40368 46572
rect 43352 46520 43404 46572
rect 44824 46520 44876 46572
rect 45836 46563 45888 46572
rect 45836 46529 45845 46563
rect 45845 46529 45879 46563
rect 45879 46529 45888 46563
rect 45836 46520 45888 46529
rect 39488 46495 39540 46504
rect 39488 46461 39497 46495
rect 39497 46461 39531 46495
rect 39531 46461 39540 46495
rect 39488 46452 39540 46461
rect 40684 46495 40736 46504
rect 40684 46461 40693 46495
rect 40693 46461 40727 46495
rect 40727 46461 40736 46495
rect 40684 46452 40736 46461
rect 41512 46452 41564 46504
rect 37372 46384 37424 46436
rect 35624 46316 35676 46368
rect 38936 46316 38988 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 11704 46112 11756 46164
rect 17592 46112 17644 46164
rect 18696 46155 18748 46164
rect 16120 46044 16172 46096
rect 18696 46121 18705 46155
rect 18705 46121 18739 46155
rect 18739 46121 18748 46155
rect 18696 46112 18748 46121
rect 24860 46112 24912 46164
rect 27068 46112 27120 46164
rect 27712 46112 27764 46164
rect 29644 46112 29696 46164
rect 31300 46112 31352 46164
rect 17408 45951 17460 45960
rect 17408 45917 17417 45951
rect 17417 45917 17451 45951
rect 17451 45917 17460 45951
rect 17408 45908 17460 45917
rect 19340 45976 19392 46028
rect 21180 46044 21232 46096
rect 24768 46044 24820 46096
rect 24308 45976 24360 46028
rect 12808 45840 12860 45892
rect 19800 45908 19852 45960
rect 19892 45908 19944 45960
rect 21732 45951 21784 45960
rect 21088 45840 21140 45892
rect 19432 45772 19484 45824
rect 19892 45772 19944 45824
rect 20628 45772 20680 45824
rect 21732 45917 21741 45951
rect 21741 45917 21775 45951
rect 21775 45917 21784 45951
rect 21732 45908 21784 45917
rect 21824 45951 21876 45960
rect 21824 45917 21837 45951
rect 21837 45917 21871 45951
rect 21871 45917 21876 45951
rect 21824 45908 21876 45917
rect 22744 45908 22796 45960
rect 23204 45908 23256 45960
rect 26148 45976 26200 46028
rect 23112 45840 23164 45892
rect 24584 45883 24636 45892
rect 24584 45849 24593 45883
rect 24593 45849 24627 45883
rect 24627 45849 24636 45883
rect 24584 45840 24636 45849
rect 26056 45908 26108 45960
rect 26240 45951 26292 45960
rect 26240 45917 26249 45951
rect 26249 45917 26283 45951
rect 26283 45917 26292 45951
rect 26240 45908 26292 45917
rect 26332 45951 26384 45960
rect 26332 45917 26341 45951
rect 26341 45917 26375 45951
rect 26375 45917 26384 45951
rect 26332 45908 26384 45917
rect 26424 45840 26476 45892
rect 26976 45951 27028 45960
rect 26976 45917 26985 45951
rect 26985 45917 27019 45951
rect 27019 45917 27028 45951
rect 29368 46044 29420 46096
rect 30932 46044 30984 46096
rect 33232 46112 33284 46164
rect 34336 46112 34388 46164
rect 35716 46112 35768 46164
rect 36360 46155 36412 46164
rect 36360 46121 36369 46155
rect 36369 46121 36403 46155
rect 36403 46121 36412 46155
rect 36360 46112 36412 46121
rect 39304 46112 39356 46164
rect 42616 46112 42668 46164
rect 44272 46155 44324 46164
rect 44272 46121 44281 46155
rect 44281 46121 44315 46155
rect 44315 46121 44324 46155
rect 44272 46112 44324 46121
rect 27896 45976 27948 46028
rect 28908 45951 28960 45960
rect 26976 45908 27028 45917
rect 28908 45917 28917 45951
rect 28917 45917 28951 45951
rect 28951 45917 28960 45951
rect 28908 45908 28960 45917
rect 27620 45840 27672 45892
rect 29000 45883 29052 45892
rect 29000 45849 29009 45883
rect 29009 45849 29043 45883
rect 29043 45849 29052 45883
rect 29000 45840 29052 45849
rect 29368 45908 29420 45960
rect 29828 45908 29880 45960
rect 30288 45908 30340 45960
rect 33140 45976 33192 46028
rect 33508 45976 33560 46028
rect 41144 46044 41196 46096
rect 32036 45951 32088 45960
rect 32036 45917 32045 45951
rect 32045 45917 32079 45951
rect 32079 45917 32088 45951
rect 32036 45908 32088 45917
rect 33416 45908 33468 45960
rect 33692 45908 33744 45960
rect 33876 45951 33928 45960
rect 33876 45917 33885 45951
rect 33885 45917 33919 45951
rect 33919 45917 33928 45951
rect 33876 45908 33928 45917
rect 30196 45840 30248 45892
rect 31944 45840 31996 45892
rect 34060 45883 34112 45892
rect 34060 45849 34069 45883
rect 34069 45849 34103 45883
rect 34103 45849 34112 45883
rect 34060 45840 34112 45849
rect 25412 45772 25464 45824
rect 27804 45772 27856 45824
rect 31484 45772 31536 45824
rect 36912 45951 36964 45960
rect 36912 45917 36921 45951
rect 36921 45917 36955 45951
rect 36955 45917 36964 45951
rect 36912 45908 36964 45917
rect 37556 45976 37608 46028
rect 38476 45976 38528 46028
rect 39488 45976 39540 46028
rect 40592 46019 40644 46028
rect 40592 45985 40601 46019
rect 40601 45985 40635 46019
rect 40635 45985 40644 46019
rect 40592 45976 40644 45985
rect 42248 45976 42300 46028
rect 37648 45908 37700 45960
rect 38568 45908 38620 45960
rect 39120 45951 39172 45960
rect 39120 45917 39129 45951
rect 39129 45917 39163 45951
rect 39163 45917 39172 45951
rect 39120 45908 39172 45917
rect 39580 45908 39632 45960
rect 34428 45840 34480 45892
rect 38108 45840 38160 45892
rect 38200 45840 38252 45892
rect 40132 45840 40184 45892
rect 40776 45908 40828 45960
rect 41236 45951 41288 45960
rect 41236 45917 41245 45951
rect 41245 45917 41279 45951
rect 41279 45917 41288 45951
rect 41236 45908 41288 45917
rect 42248 45840 42300 45892
rect 41420 45772 41472 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 17132 45568 17184 45620
rect 19340 45568 19392 45620
rect 20536 45568 20588 45620
rect 20628 45568 20680 45620
rect 17960 45432 18012 45484
rect 18788 45475 18840 45484
rect 18788 45441 18797 45475
rect 18797 45441 18831 45475
rect 18831 45441 18840 45475
rect 18788 45432 18840 45441
rect 18972 45475 19024 45484
rect 18972 45441 18981 45475
rect 18981 45441 19015 45475
rect 19015 45441 19024 45475
rect 18972 45432 19024 45441
rect 20904 45475 20956 45484
rect 20904 45441 20913 45475
rect 20913 45441 20947 45475
rect 20947 45441 20956 45475
rect 20904 45432 20956 45441
rect 20996 45432 21048 45484
rect 23848 45568 23900 45620
rect 24308 45568 24360 45620
rect 27528 45568 27580 45620
rect 29276 45568 29328 45620
rect 23480 45500 23532 45552
rect 24584 45500 24636 45552
rect 25136 45500 25188 45552
rect 25320 45500 25372 45552
rect 4620 45364 4672 45416
rect 20168 45364 20220 45416
rect 20628 45296 20680 45348
rect 23204 45475 23256 45484
rect 23204 45441 23213 45475
rect 23213 45441 23247 45475
rect 23247 45441 23256 45475
rect 23204 45432 23256 45441
rect 25412 45432 25464 45484
rect 26056 45475 26108 45484
rect 23020 45364 23072 45416
rect 23112 45407 23164 45416
rect 23112 45373 23121 45407
rect 23121 45373 23155 45407
rect 23155 45373 23164 45407
rect 23112 45364 23164 45373
rect 26056 45441 26065 45475
rect 26065 45441 26099 45475
rect 26099 45441 26108 45475
rect 26056 45432 26108 45441
rect 26148 45432 26200 45484
rect 25504 45296 25556 45348
rect 26424 45364 26476 45416
rect 28448 45364 28500 45416
rect 28908 45432 28960 45484
rect 29000 45364 29052 45416
rect 29920 45432 29972 45484
rect 30012 45432 30064 45484
rect 31024 45475 31076 45484
rect 31024 45441 31033 45475
rect 31033 45441 31067 45475
rect 31067 45441 31076 45475
rect 31024 45432 31076 45441
rect 36268 45568 36320 45620
rect 40592 45568 40644 45620
rect 41236 45568 41288 45620
rect 43904 45568 43956 45620
rect 45192 45568 45244 45620
rect 34796 45500 34848 45552
rect 33048 45432 33100 45484
rect 33416 45432 33468 45484
rect 35624 45500 35676 45552
rect 36636 45500 36688 45552
rect 41788 45500 41840 45552
rect 29736 45364 29788 45416
rect 34060 45407 34112 45416
rect 34060 45373 34069 45407
rect 34069 45373 34103 45407
rect 34103 45373 34112 45407
rect 34060 45364 34112 45373
rect 36728 45475 36780 45484
rect 35532 45364 35584 45416
rect 35716 45364 35768 45416
rect 36268 45407 36320 45416
rect 36268 45373 36277 45407
rect 36277 45373 36311 45407
rect 36311 45373 36320 45407
rect 36268 45364 36320 45373
rect 26332 45296 26384 45348
rect 24216 45228 24268 45280
rect 25228 45228 25280 45280
rect 26608 45296 26660 45348
rect 27988 45339 28040 45348
rect 27988 45305 27997 45339
rect 27997 45305 28031 45339
rect 28031 45305 28040 45339
rect 27988 45296 28040 45305
rect 30380 45296 30432 45348
rect 36728 45441 36737 45475
rect 36737 45441 36771 45475
rect 36771 45441 36780 45475
rect 36728 45432 36780 45441
rect 38108 45475 38160 45484
rect 38108 45441 38117 45475
rect 38117 45441 38151 45475
rect 38151 45441 38160 45475
rect 38108 45432 38160 45441
rect 38660 45432 38712 45484
rect 39120 45475 39172 45484
rect 39120 45441 39129 45475
rect 39129 45441 39163 45475
rect 39163 45441 39172 45475
rect 39120 45432 39172 45441
rect 40316 45475 40368 45484
rect 40316 45441 40325 45475
rect 40325 45441 40359 45475
rect 40359 45441 40368 45475
rect 40316 45432 40368 45441
rect 40776 45475 40828 45484
rect 40776 45441 40785 45475
rect 40785 45441 40819 45475
rect 40819 45441 40828 45475
rect 40776 45432 40828 45441
rect 41512 45475 41564 45484
rect 41512 45441 41521 45475
rect 41521 45441 41555 45475
rect 41555 45441 41564 45475
rect 41512 45432 41564 45441
rect 42616 45475 42668 45484
rect 42616 45441 42625 45475
rect 42625 45441 42659 45475
rect 42659 45441 42668 45475
rect 42616 45432 42668 45441
rect 37188 45364 37240 45416
rect 37648 45364 37700 45416
rect 38200 45364 38252 45416
rect 38568 45407 38620 45416
rect 38568 45373 38577 45407
rect 38577 45373 38611 45407
rect 38611 45373 38620 45407
rect 38568 45364 38620 45373
rect 37372 45296 37424 45348
rect 37556 45296 37608 45348
rect 38292 45296 38344 45348
rect 27252 45271 27304 45280
rect 27252 45237 27261 45271
rect 27261 45237 27295 45271
rect 27295 45237 27304 45271
rect 27252 45228 27304 45237
rect 27804 45228 27856 45280
rect 29552 45228 29604 45280
rect 37648 45228 37700 45280
rect 40408 45364 40460 45416
rect 40592 45407 40644 45416
rect 40592 45373 40601 45407
rect 40601 45373 40635 45407
rect 40635 45373 40644 45407
rect 40592 45364 40644 45373
rect 39856 45339 39908 45348
rect 39856 45305 39865 45339
rect 39865 45305 39899 45339
rect 39899 45305 39908 45339
rect 39856 45296 39908 45305
rect 39304 45271 39356 45280
rect 39304 45237 39313 45271
rect 39313 45237 39347 45271
rect 39347 45237 39356 45271
rect 43260 45364 43312 45416
rect 39304 45228 39356 45237
rect 42708 45228 42760 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 18328 45067 18380 45076
rect 18328 45033 18337 45067
rect 18337 45033 18371 45067
rect 18371 45033 18380 45067
rect 18328 45024 18380 45033
rect 24952 45024 25004 45076
rect 25504 45024 25556 45076
rect 34152 45067 34204 45076
rect 23112 44956 23164 45008
rect 25596 44956 25648 45008
rect 26056 44956 26108 45008
rect 29736 44956 29788 45008
rect 34152 45033 34161 45067
rect 34161 45033 34195 45067
rect 34195 45033 34204 45067
rect 34152 45024 34204 45033
rect 39948 45024 40000 45076
rect 42248 45067 42300 45076
rect 42248 45033 42257 45067
rect 42257 45033 42291 45067
rect 42291 45033 42300 45067
rect 42248 45024 42300 45033
rect 20904 44888 20956 44940
rect 18144 44863 18196 44872
rect 18144 44829 18153 44863
rect 18153 44829 18187 44863
rect 18187 44829 18196 44863
rect 18144 44820 18196 44829
rect 19984 44863 20036 44872
rect 19984 44829 19993 44863
rect 19993 44829 20027 44863
rect 20027 44829 20036 44863
rect 19984 44820 20036 44829
rect 20996 44820 21048 44872
rect 22008 44863 22060 44872
rect 22008 44829 22017 44863
rect 22017 44829 22051 44863
rect 22051 44829 22060 44863
rect 22008 44820 22060 44829
rect 23020 44820 23072 44872
rect 22192 44795 22244 44804
rect 22192 44761 22201 44795
rect 22201 44761 22235 44795
rect 22235 44761 22244 44795
rect 22192 44752 22244 44761
rect 24124 44888 24176 44940
rect 25412 44931 25464 44940
rect 25412 44897 25421 44931
rect 25421 44897 25455 44931
rect 25455 44897 25464 44931
rect 25412 44888 25464 44897
rect 23480 44820 23532 44872
rect 24216 44820 24268 44872
rect 25320 44820 25372 44872
rect 25964 44863 26016 44872
rect 25964 44829 25973 44863
rect 25973 44829 26007 44863
rect 26007 44829 26016 44863
rect 25964 44820 26016 44829
rect 26240 44863 26292 44872
rect 26240 44829 26249 44863
rect 26249 44829 26283 44863
rect 26283 44829 26292 44863
rect 26240 44820 26292 44829
rect 26424 44863 26476 44872
rect 26424 44829 26433 44863
rect 26433 44829 26467 44863
rect 26467 44829 26476 44863
rect 26424 44820 26476 44829
rect 27620 44863 27672 44872
rect 27620 44829 27629 44863
rect 27629 44829 27663 44863
rect 27663 44829 27672 44863
rect 27620 44820 27672 44829
rect 27160 44795 27212 44804
rect 18788 44684 18840 44736
rect 21916 44727 21968 44736
rect 21916 44693 21925 44727
rect 21925 44693 21959 44727
rect 21959 44693 21968 44727
rect 21916 44684 21968 44693
rect 22376 44684 22428 44736
rect 24308 44684 24360 44736
rect 27160 44761 27169 44795
rect 27169 44761 27203 44795
rect 27203 44761 27212 44795
rect 27160 44752 27212 44761
rect 29644 44888 29696 44940
rect 30288 44888 30340 44940
rect 34980 44956 35032 45008
rect 35348 44956 35400 45008
rect 27988 44863 28040 44872
rect 27988 44829 27997 44863
rect 27997 44829 28031 44863
rect 28031 44829 28040 44863
rect 27988 44820 28040 44829
rect 29552 44820 29604 44872
rect 33416 44888 33468 44940
rect 31944 44863 31996 44872
rect 31944 44829 31953 44863
rect 31953 44829 31987 44863
rect 31987 44829 31996 44863
rect 31944 44820 31996 44829
rect 32036 44863 32088 44872
rect 32036 44829 32045 44863
rect 32045 44829 32079 44863
rect 32079 44829 32088 44863
rect 32312 44863 32364 44872
rect 32036 44820 32088 44829
rect 32312 44829 32321 44863
rect 32321 44829 32355 44863
rect 32355 44829 32364 44863
rect 32312 44820 32364 44829
rect 34060 44888 34112 44940
rect 36268 44888 36320 44940
rect 33968 44820 34020 44872
rect 35532 44863 35584 44872
rect 33140 44795 33192 44804
rect 28172 44684 28224 44736
rect 33140 44761 33149 44795
rect 33149 44761 33183 44795
rect 33183 44761 33192 44795
rect 33140 44752 33192 44761
rect 34612 44684 34664 44736
rect 35532 44829 35541 44863
rect 35541 44829 35575 44863
rect 35575 44829 35584 44863
rect 35532 44820 35584 44829
rect 35716 44863 35768 44872
rect 35716 44829 35725 44863
rect 35725 44829 35759 44863
rect 35759 44829 35768 44863
rect 35716 44820 35768 44829
rect 37372 44820 37424 44872
rect 37556 44820 37608 44872
rect 38660 44863 38712 44872
rect 36452 44795 36504 44804
rect 36452 44761 36461 44795
rect 36461 44761 36495 44795
rect 36495 44761 36504 44795
rect 36452 44752 36504 44761
rect 38660 44829 38669 44863
rect 38669 44829 38703 44863
rect 38703 44829 38712 44863
rect 38660 44820 38712 44829
rect 39488 44888 39540 44940
rect 40316 44888 40368 44940
rect 41420 44888 41472 44940
rect 42708 44931 42760 44940
rect 39304 44863 39356 44872
rect 39304 44829 39313 44863
rect 39313 44829 39347 44863
rect 39347 44829 39356 44863
rect 39304 44820 39356 44829
rect 41328 44820 41380 44872
rect 42708 44897 42717 44931
rect 42717 44897 42751 44931
rect 42751 44897 42760 44931
rect 42708 44888 42760 44897
rect 40776 44752 40828 44804
rect 36176 44684 36228 44736
rect 37188 44684 37240 44736
rect 40224 44684 40276 44736
rect 43260 44727 43312 44736
rect 43260 44693 43269 44727
rect 43269 44693 43303 44727
rect 43303 44693 43312 44727
rect 43260 44684 43312 44693
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 18972 44480 19024 44532
rect 20536 44480 20588 44532
rect 22008 44480 22060 44532
rect 22376 44480 22428 44532
rect 18052 44412 18104 44464
rect 19064 44387 19116 44396
rect 19064 44353 19073 44387
rect 19073 44353 19107 44387
rect 19107 44353 19116 44387
rect 19064 44344 19116 44353
rect 19984 44344 20036 44396
rect 20536 44387 20588 44396
rect 20536 44353 20545 44387
rect 20545 44353 20579 44387
rect 20579 44353 20588 44387
rect 20536 44344 20588 44353
rect 21088 44387 21140 44396
rect 21088 44353 21097 44387
rect 21097 44353 21131 44387
rect 21131 44353 21140 44387
rect 21088 44344 21140 44353
rect 21916 44412 21968 44464
rect 22652 44412 22704 44464
rect 20720 44276 20772 44328
rect 23112 44480 23164 44532
rect 24216 44480 24268 44532
rect 26332 44523 26384 44532
rect 22836 44455 22888 44464
rect 22836 44421 22845 44455
rect 22845 44421 22879 44455
rect 22879 44421 22888 44455
rect 22836 44412 22888 44421
rect 23020 44412 23072 44464
rect 26332 44489 26341 44523
rect 26341 44489 26375 44523
rect 26375 44489 26384 44523
rect 26332 44480 26384 44489
rect 27804 44480 27856 44532
rect 22928 44387 22980 44396
rect 22928 44353 22937 44387
rect 22937 44353 22971 44387
rect 22971 44353 22980 44387
rect 22928 44344 22980 44353
rect 24308 44387 24360 44396
rect 24308 44353 24317 44387
rect 24317 44353 24351 44387
rect 24351 44353 24360 44387
rect 24308 44344 24360 44353
rect 24768 44387 24820 44396
rect 24768 44353 24777 44387
rect 24777 44353 24811 44387
rect 24811 44353 24820 44387
rect 24768 44344 24820 44353
rect 25228 44387 25280 44396
rect 25228 44353 25237 44387
rect 25237 44353 25271 44387
rect 25271 44353 25280 44387
rect 25228 44344 25280 44353
rect 26056 44344 26108 44396
rect 27988 44412 28040 44464
rect 27620 44344 27672 44396
rect 23112 44319 23164 44328
rect 23112 44285 23121 44319
rect 23121 44285 23155 44319
rect 23155 44285 23164 44319
rect 23112 44276 23164 44285
rect 27344 44276 27396 44328
rect 39856 44480 39908 44532
rect 41328 44480 41380 44532
rect 42248 44480 42300 44532
rect 29092 44412 29144 44464
rect 33416 44455 33468 44464
rect 28448 44344 28500 44396
rect 29828 44387 29880 44396
rect 29000 44319 29052 44328
rect 29000 44285 29009 44319
rect 29009 44285 29043 44319
rect 29043 44285 29052 44319
rect 29000 44276 29052 44285
rect 29828 44353 29837 44387
rect 29837 44353 29871 44387
rect 29871 44353 29880 44387
rect 29828 44344 29880 44353
rect 33416 44421 33425 44455
rect 33425 44421 33459 44455
rect 33459 44421 33468 44455
rect 33416 44412 33468 44421
rect 34428 44412 34480 44464
rect 34980 44455 35032 44464
rect 34980 44421 34989 44455
rect 34989 44421 35023 44455
rect 35023 44421 35032 44455
rect 34980 44412 35032 44421
rect 29736 44276 29788 44328
rect 28172 44208 28224 44260
rect 31576 44208 31628 44260
rect 31944 44344 31996 44396
rect 34336 44387 34388 44396
rect 34336 44353 34345 44387
rect 34345 44353 34379 44387
rect 34379 44353 34388 44387
rect 34336 44344 34388 44353
rect 34612 44344 34664 44396
rect 35624 44387 35676 44396
rect 35624 44353 35633 44387
rect 35633 44353 35667 44387
rect 35667 44353 35676 44387
rect 35624 44344 35676 44353
rect 36176 44387 36228 44396
rect 36176 44353 36185 44387
rect 36185 44353 36219 44387
rect 36219 44353 36228 44387
rect 36176 44344 36228 44353
rect 31852 44276 31904 44328
rect 33140 44276 33192 44328
rect 33692 44276 33744 44328
rect 34796 44276 34848 44328
rect 35716 44276 35768 44328
rect 38292 44387 38344 44396
rect 36360 44319 36412 44328
rect 36360 44285 36369 44319
rect 36369 44285 36403 44319
rect 36403 44285 36412 44319
rect 36360 44276 36412 44285
rect 32036 44140 32088 44192
rect 38292 44353 38301 44387
rect 38301 44353 38335 44387
rect 38335 44353 38344 44387
rect 38292 44344 38344 44353
rect 38476 44276 38528 44328
rect 40408 44412 40460 44464
rect 40592 44344 40644 44396
rect 40776 44344 40828 44396
rect 39948 44276 40000 44328
rect 34152 44140 34204 44192
rect 34428 44140 34480 44192
rect 41880 44208 41932 44260
rect 39396 44183 39448 44192
rect 39396 44149 39405 44183
rect 39405 44149 39439 44183
rect 39439 44149 39448 44183
rect 39396 44140 39448 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 21732 43936 21784 43988
rect 20536 43868 20588 43920
rect 24400 43936 24452 43988
rect 28264 43936 28316 43988
rect 30104 43979 30156 43988
rect 30104 43945 30113 43979
rect 30113 43945 30147 43979
rect 30147 43945 30156 43979
rect 30104 43936 30156 43945
rect 31116 43979 31168 43988
rect 31116 43945 31125 43979
rect 31125 43945 31159 43979
rect 31159 43945 31168 43979
rect 31116 43936 31168 43945
rect 31760 43936 31812 43988
rect 32312 43936 32364 43988
rect 37280 43979 37332 43988
rect 37280 43945 37289 43979
rect 37289 43945 37323 43979
rect 37323 43945 37332 43979
rect 37280 43936 37332 43945
rect 38476 43936 38528 43988
rect 40592 43979 40644 43988
rect 40592 43945 40601 43979
rect 40601 43945 40635 43979
rect 40635 43945 40644 43979
rect 40592 43936 40644 43945
rect 43260 43936 43312 43988
rect 20168 43843 20220 43852
rect 20168 43809 20177 43843
rect 20177 43809 20211 43843
rect 20211 43809 20220 43843
rect 20168 43800 20220 43809
rect 20536 43775 20588 43784
rect 20536 43741 20545 43775
rect 20545 43741 20579 43775
rect 20579 43741 20588 43775
rect 20536 43732 20588 43741
rect 20720 43775 20772 43784
rect 20720 43741 20729 43775
rect 20729 43741 20763 43775
rect 20763 43741 20772 43775
rect 20720 43732 20772 43741
rect 21916 43800 21968 43852
rect 27252 43868 27304 43920
rect 30564 43868 30616 43920
rect 22744 43732 22796 43784
rect 33692 43843 33744 43852
rect 33692 43809 33701 43843
rect 33701 43809 33735 43843
rect 33735 43809 33744 43843
rect 33692 43800 33744 43809
rect 38108 43800 38160 43852
rect 24768 43732 24820 43784
rect 23112 43664 23164 43716
rect 23296 43707 23348 43716
rect 23296 43673 23305 43707
rect 23305 43673 23339 43707
rect 23339 43673 23348 43707
rect 23296 43664 23348 43673
rect 23388 43664 23440 43716
rect 27344 43732 27396 43784
rect 27620 43775 27672 43784
rect 27620 43741 27629 43775
rect 27629 43741 27663 43775
rect 27663 43741 27672 43775
rect 27620 43732 27672 43741
rect 27804 43775 27856 43784
rect 27804 43741 27813 43775
rect 27813 43741 27847 43775
rect 27847 43741 27856 43775
rect 27804 43732 27856 43741
rect 28080 43775 28132 43784
rect 28080 43741 28089 43775
rect 28089 43741 28123 43775
rect 28123 43741 28132 43775
rect 28080 43732 28132 43741
rect 28172 43732 28224 43784
rect 31852 43732 31904 43784
rect 32772 43732 32824 43784
rect 33784 43775 33836 43784
rect 33784 43741 33793 43775
rect 33793 43741 33827 43775
rect 33827 43741 33836 43775
rect 33784 43732 33836 43741
rect 34152 43775 34204 43784
rect 34152 43741 34161 43775
rect 34161 43741 34195 43775
rect 34195 43741 34204 43775
rect 34152 43732 34204 43741
rect 34520 43732 34572 43784
rect 34796 43732 34848 43784
rect 27988 43664 28040 43716
rect 34428 43664 34480 43716
rect 38568 43775 38620 43784
rect 35532 43664 35584 43716
rect 20628 43596 20680 43648
rect 21180 43596 21232 43648
rect 23020 43639 23072 43648
rect 23020 43605 23029 43639
rect 23029 43605 23063 43639
rect 23063 43605 23072 43639
rect 23020 43596 23072 43605
rect 34612 43596 34664 43648
rect 38568 43741 38577 43775
rect 38577 43741 38611 43775
rect 38611 43741 38620 43775
rect 38568 43732 38620 43741
rect 38660 43775 38712 43784
rect 38660 43741 38669 43775
rect 38669 43741 38703 43775
rect 38703 43741 38712 43775
rect 38660 43732 38712 43741
rect 41144 43639 41196 43648
rect 41144 43605 41153 43639
rect 41153 43605 41187 43639
rect 41187 43605 41196 43639
rect 41144 43596 41196 43605
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 28172 43435 28224 43444
rect 28172 43401 28181 43435
rect 28181 43401 28215 43435
rect 28215 43401 28224 43435
rect 28172 43392 28224 43401
rect 23112 43324 23164 43376
rect 21272 43299 21324 43308
rect 21272 43265 21281 43299
rect 21281 43265 21315 43299
rect 21315 43265 21324 43299
rect 21272 43256 21324 43265
rect 22192 43256 22244 43308
rect 23388 43256 23440 43308
rect 23756 43256 23808 43308
rect 24032 43299 24084 43308
rect 24032 43265 24041 43299
rect 24041 43265 24075 43299
rect 24075 43265 24084 43299
rect 24032 43256 24084 43265
rect 24584 43324 24636 43376
rect 25228 43256 25280 43308
rect 26056 43256 26108 43308
rect 27620 43324 27672 43376
rect 22008 43231 22060 43240
rect 22008 43197 22017 43231
rect 22017 43197 22051 43231
rect 22051 43197 22060 43231
rect 22008 43188 22060 43197
rect 23296 43188 23348 43240
rect 27160 43256 27212 43308
rect 27804 43256 27856 43308
rect 28540 43256 28592 43308
rect 30380 43324 30432 43376
rect 32772 43367 32824 43376
rect 32772 43333 32781 43367
rect 32781 43333 32815 43367
rect 32815 43333 32824 43367
rect 32772 43324 32824 43333
rect 27620 43188 27672 43240
rect 27988 43188 28040 43240
rect 23664 43120 23716 43172
rect 27252 43120 27304 43172
rect 30012 43299 30064 43308
rect 30012 43265 30021 43299
rect 30021 43265 30055 43299
rect 30055 43265 30064 43299
rect 30012 43256 30064 43265
rect 30564 43256 30616 43308
rect 34152 43324 34204 43376
rect 34244 43299 34296 43308
rect 29736 43231 29788 43240
rect 29736 43197 29745 43231
rect 29745 43197 29779 43231
rect 29779 43197 29788 43231
rect 29736 43188 29788 43197
rect 31300 43120 31352 43172
rect 34244 43265 34253 43299
rect 34253 43265 34287 43299
rect 34287 43265 34296 43299
rect 34244 43256 34296 43265
rect 36728 43324 36780 43376
rect 37464 43324 37516 43376
rect 36452 43256 36504 43308
rect 39396 43299 39448 43308
rect 39396 43265 39405 43299
rect 39405 43265 39439 43299
rect 39439 43265 39448 43299
rect 39396 43256 39448 43265
rect 39948 43299 40000 43308
rect 39948 43265 39957 43299
rect 39957 43265 39991 43299
rect 39991 43265 40000 43299
rect 39948 43256 40000 43265
rect 34520 43188 34572 43240
rect 33784 43120 33836 43172
rect 34612 43052 34664 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 23204 42891 23256 42900
rect 23204 42857 23213 42891
rect 23213 42857 23247 42891
rect 23247 42857 23256 42891
rect 23204 42848 23256 42857
rect 25228 42848 25280 42900
rect 22652 42687 22704 42696
rect 22652 42653 22661 42687
rect 22661 42653 22695 42687
rect 22695 42653 22704 42687
rect 22652 42644 22704 42653
rect 23020 42687 23072 42696
rect 23020 42653 23029 42687
rect 23029 42653 23063 42687
rect 23063 42653 23072 42687
rect 23020 42644 23072 42653
rect 25412 42687 25464 42696
rect 25412 42653 25421 42687
rect 25421 42653 25455 42687
rect 25455 42653 25464 42687
rect 25412 42644 25464 42653
rect 26240 42848 26292 42900
rect 29644 42780 29696 42832
rect 30012 42780 30064 42832
rect 28080 42712 28132 42764
rect 29736 42712 29788 42764
rect 33140 42755 33192 42764
rect 33140 42721 33149 42755
rect 33149 42721 33183 42755
rect 33183 42721 33192 42755
rect 33140 42712 33192 42721
rect 33784 42755 33836 42764
rect 33784 42721 33793 42755
rect 33793 42721 33827 42755
rect 33827 42721 33836 42755
rect 33784 42712 33836 42721
rect 27620 42644 27672 42696
rect 27988 42687 28040 42696
rect 27988 42653 27997 42687
rect 27997 42653 28031 42687
rect 28031 42653 28040 42687
rect 27988 42644 28040 42653
rect 28172 42644 28224 42696
rect 23756 42576 23808 42628
rect 27160 42576 27212 42628
rect 22928 42508 22980 42560
rect 30380 42644 30432 42696
rect 32404 42687 32456 42696
rect 32404 42653 32413 42687
rect 32413 42653 32447 42687
rect 32447 42653 32456 42687
rect 32404 42644 32456 42653
rect 33416 42644 33468 42696
rect 34612 42712 34664 42764
rect 34704 42712 34756 42764
rect 35440 42712 35492 42764
rect 37556 42712 37608 42764
rect 40132 42712 40184 42764
rect 41144 42712 41196 42764
rect 34336 42687 34388 42696
rect 34336 42653 34345 42687
rect 34345 42653 34379 42687
rect 34379 42653 34388 42687
rect 34336 42644 34388 42653
rect 37188 42644 37240 42696
rect 29460 42576 29512 42628
rect 30196 42576 30248 42628
rect 30656 42508 30708 42560
rect 36912 42551 36964 42560
rect 36912 42517 36921 42551
rect 36921 42517 36955 42551
rect 36955 42517 36964 42551
rect 36912 42508 36964 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 22652 42304 22704 42356
rect 26240 42347 26292 42356
rect 23756 42211 23808 42220
rect 23756 42177 23765 42211
rect 23765 42177 23799 42211
rect 23799 42177 23808 42211
rect 23756 42168 23808 42177
rect 24032 42168 24084 42220
rect 26240 42313 26249 42347
rect 26249 42313 26283 42347
rect 26283 42313 26292 42347
rect 26240 42304 26292 42313
rect 25412 42236 25464 42288
rect 30564 42304 30616 42356
rect 30656 42347 30708 42356
rect 30656 42313 30665 42347
rect 30665 42313 30699 42347
rect 30699 42313 30708 42347
rect 30656 42304 30708 42313
rect 31024 42304 31076 42356
rect 33968 42304 34020 42356
rect 34336 42304 34388 42356
rect 36912 42304 36964 42356
rect 38108 42347 38160 42356
rect 38108 42313 38117 42347
rect 38117 42313 38151 42347
rect 38151 42313 38160 42347
rect 38108 42304 38160 42313
rect 36728 42279 36780 42288
rect 36728 42245 36737 42279
rect 36737 42245 36771 42279
rect 36771 42245 36780 42279
rect 36728 42236 36780 42245
rect 24584 42143 24636 42152
rect 24584 42109 24593 42143
rect 24593 42109 24627 42143
rect 24627 42109 24636 42143
rect 24584 42100 24636 42109
rect 29460 42211 29512 42220
rect 29460 42177 29469 42211
rect 29469 42177 29503 42211
rect 29503 42177 29512 42211
rect 29460 42168 29512 42177
rect 30656 42168 30708 42220
rect 32220 42168 32272 42220
rect 22008 41964 22060 42016
rect 22744 41964 22796 42016
rect 26608 41964 26660 42016
rect 35532 42007 35584 42016
rect 35532 41973 35541 42007
rect 35541 41973 35575 42007
rect 35575 41973 35584 42007
rect 35532 41964 35584 41973
rect 37188 41964 37240 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 24768 41760 24820 41812
rect 28172 41760 28224 41812
rect 31300 41803 31352 41812
rect 31300 41769 31309 41803
rect 31309 41769 31343 41803
rect 31343 41769 31352 41803
rect 31300 41760 31352 41769
rect 33968 41760 34020 41812
rect 33140 41692 33192 41744
rect 35532 41692 35584 41744
rect 26240 41556 26292 41608
rect 26608 41599 26660 41608
rect 26608 41565 26617 41599
rect 26617 41565 26651 41599
rect 26651 41565 26660 41599
rect 26608 41556 26660 41565
rect 27620 41488 27672 41540
rect 30472 41488 30524 41540
rect 30840 41531 30892 41540
rect 30840 41497 30849 41531
rect 30849 41497 30883 41531
rect 30883 41497 30892 41531
rect 30840 41488 30892 41497
rect 27344 41420 27396 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 22744 41216 22796 41268
rect 26240 41216 26292 41268
rect 26516 41259 26568 41268
rect 26516 41225 26525 41259
rect 26525 41225 26559 41259
rect 26559 41225 26568 41259
rect 26516 41216 26568 41225
rect 27344 41216 27396 41268
rect 28540 41259 28592 41268
rect 28540 41225 28549 41259
rect 28549 41225 28583 41259
rect 28583 41225 28592 41259
rect 28540 41216 28592 41225
rect 32404 41216 32456 41268
rect 25964 41148 26016 41200
rect 30196 41148 30248 41200
rect 26240 41080 26292 41132
rect 29644 40919 29696 40928
rect 29644 40885 29653 40919
rect 29653 40885 29687 40919
rect 29687 40885 29696 40919
rect 29644 40876 29696 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 29644 40672 29696 40724
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 23020 7828 23072 7880
rect 24032 7871 24084 7880
rect 24032 7837 24041 7871
rect 24041 7837 24075 7871
rect 24075 7837 24084 7871
rect 24032 7828 24084 7837
rect 24952 7828 25004 7880
rect 26056 7871 26108 7880
rect 26056 7837 26065 7871
rect 26065 7837 26099 7871
rect 26099 7837 26108 7871
rect 26056 7828 26108 7837
rect 26148 7760 26200 7812
rect 25412 7735 25464 7744
rect 25412 7701 25421 7735
rect 25421 7701 25455 7735
rect 25455 7701 25464 7735
rect 25412 7692 25464 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 21272 7531 21324 7540
rect 21272 7497 21281 7531
rect 21281 7497 21315 7531
rect 21315 7497 21324 7531
rect 21272 7488 21324 7497
rect 24860 7463 24912 7472
rect 24860 7429 24869 7463
rect 24869 7429 24903 7463
rect 24903 7429 24912 7463
rect 24860 7420 24912 7429
rect 24952 7463 25004 7472
rect 24952 7429 24961 7463
rect 24961 7429 24995 7463
rect 24995 7429 25004 7463
rect 25688 7463 25740 7472
rect 24952 7420 25004 7429
rect 25688 7429 25697 7463
rect 25697 7429 25731 7463
rect 25731 7429 25740 7463
rect 25688 7420 25740 7429
rect 22100 7352 22152 7404
rect 25228 7284 25280 7336
rect 26056 7284 26108 7336
rect 26608 7327 26660 7336
rect 26608 7293 26617 7327
rect 26617 7293 26651 7327
rect 26651 7293 26660 7327
rect 26608 7284 26660 7293
rect 22468 7148 22520 7200
rect 23112 7148 23164 7200
rect 26240 7148 26292 7200
rect 27712 7148 27764 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 24860 6987 24912 6996
rect 24860 6953 24869 6987
rect 24869 6953 24903 6987
rect 24903 6953 24912 6987
rect 24860 6944 24912 6953
rect 25688 6987 25740 6996
rect 25688 6953 25697 6987
rect 25697 6953 25731 6987
rect 25731 6953 25740 6987
rect 25688 6944 25740 6953
rect 23020 6851 23072 6860
rect 23020 6817 23029 6851
rect 23029 6817 23063 6851
rect 23063 6817 23072 6851
rect 23020 6808 23072 6817
rect 23848 6851 23900 6860
rect 23848 6817 23857 6851
rect 23857 6817 23891 6851
rect 23891 6817 23900 6851
rect 23848 6808 23900 6817
rect 27712 6851 27764 6860
rect 27712 6817 27721 6851
rect 27721 6817 27755 6851
rect 27755 6817 27764 6851
rect 27712 6808 27764 6817
rect 27988 6851 28040 6860
rect 27988 6817 27997 6851
rect 27997 6817 28031 6851
rect 28031 6817 28040 6851
rect 27988 6808 28040 6817
rect 19340 6604 19392 6656
rect 21272 6740 21324 6792
rect 20904 6647 20956 6656
rect 20904 6613 20913 6647
rect 20913 6613 20947 6647
rect 20947 6613 20956 6647
rect 20904 6604 20956 6613
rect 21548 6604 21600 6656
rect 22100 6604 22152 6656
rect 22284 6647 22336 6656
rect 22284 6613 22293 6647
rect 22293 6613 22327 6647
rect 22327 6613 22336 6647
rect 22284 6604 22336 6613
rect 23112 6715 23164 6724
rect 23112 6681 23121 6715
rect 23121 6681 23155 6715
rect 23155 6681 23164 6715
rect 23112 6672 23164 6681
rect 23388 6672 23440 6724
rect 25412 6740 25464 6792
rect 26148 6604 26200 6656
rect 27804 6715 27856 6724
rect 27804 6681 27813 6715
rect 27813 6681 27847 6715
rect 27847 6681 27856 6715
rect 27804 6672 27856 6681
rect 29000 6604 29052 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 27804 6400 27856 6452
rect 20536 6375 20588 6384
rect 20536 6341 20545 6375
rect 20545 6341 20579 6375
rect 20579 6341 20588 6375
rect 20536 6332 20588 6341
rect 22560 6375 22612 6384
rect 22560 6341 22569 6375
rect 22569 6341 22603 6375
rect 22603 6341 22612 6375
rect 22560 6332 22612 6341
rect 24032 6375 24084 6384
rect 24032 6341 24041 6375
rect 24041 6341 24075 6375
rect 24075 6341 24084 6375
rect 24032 6332 24084 6341
rect 24124 6375 24176 6384
rect 24124 6341 24133 6375
rect 24133 6341 24167 6375
rect 24167 6341 24176 6375
rect 25688 6375 25740 6384
rect 24124 6332 24176 6341
rect 25688 6341 25697 6375
rect 25697 6341 25731 6375
rect 25731 6341 25740 6375
rect 25688 6332 25740 6341
rect 26516 6264 26568 6316
rect 21088 6239 21140 6248
rect 21088 6205 21097 6239
rect 21097 6205 21131 6239
rect 21131 6205 21140 6239
rect 21088 6196 21140 6205
rect 22468 6239 22520 6248
rect 22468 6205 22477 6239
rect 22477 6205 22511 6239
rect 22511 6205 22520 6239
rect 22468 6196 22520 6205
rect 23572 6196 23624 6248
rect 24952 6239 25004 6248
rect 24952 6205 24961 6239
rect 24961 6205 24995 6239
rect 24995 6205 25004 6239
rect 24952 6196 25004 6205
rect 26240 6196 26292 6248
rect 26332 6128 26384 6180
rect 28172 6060 28224 6112
rect 29736 6060 29788 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 20536 5856 20588 5908
rect 22560 5899 22612 5908
rect 22560 5865 22569 5899
rect 22569 5865 22603 5899
rect 22603 5865 22612 5899
rect 22560 5856 22612 5865
rect 24124 5856 24176 5908
rect 25688 5899 25740 5908
rect 25688 5865 25697 5899
rect 25697 5865 25731 5899
rect 25731 5865 25740 5899
rect 25688 5856 25740 5865
rect 26516 5856 26568 5908
rect 22284 5720 22336 5772
rect 26148 5720 26200 5772
rect 27712 5763 27764 5772
rect 20352 5652 20404 5704
rect 20904 5695 20956 5704
rect 20904 5661 20913 5695
rect 20913 5661 20947 5695
rect 20947 5661 20956 5695
rect 20904 5652 20956 5661
rect 21548 5652 21600 5704
rect 22836 5652 22888 5704
rect 23388 5652 23440 5704
rect 25412 5695 25464 5704
rect 25412 5661 25421 5695
rect 25421 5661 25455 5695
rect 25455 5661 25464 5695
rect 25412 5652 25464 5661
rect 27712 5729 27721 5763
rect 27721 5729 27755 5763
rect 27755 5729 27764 5763
rect 27712 5720 27764 5729
rect 29000 5695 29052 5704
rect 29000 5661 29009 5695
rect 29009 5661 29043 5695
rect 29043 5661 29052 5695
rect 29000 5652 29052 5661
rect 22652 5584 22704 5636
rect 24308 5584 24360 5636
rect 28172 5627 28224 5636
rect 28172 5593 28181 5627
rect 28181 5593 28215 5627
rect 28215 5593 28224 5627
rect 28172 5584 28224 5593
rect 28264 5627 28316 5636
rect 28264 5593 28273 5627
rect 28273 5593 28307 5627
rect 28307 5593 28316 5627
rect 28264 5584 28316 5593
rect 29644 5584 29696 5636
rect 20076 5559 20128 5568
rect 20076 5525 20085 5559
rect 20085 5525 20119 5559
rect 20119 5525 20128 5559
rect 20076 5516 20128 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 20076 5244 20128 5296
rect 22652 5287 22704 5296
rect 22652 5253 22661 5287
rect 22661 5253 22695 5287
rect 22695 5253 22704 5287
rect 22652 5244 22704 5253
rect 24308 5287 24360 5296
rect 24308 5253 24317 5287
rect 24317 5253 24351 5287
rect 24351 5253 24360 5287
rect 24308 5244 24360 5253
rect 29644 5287 29696 5296
rect 29644 5253 29653 5287
rect 29653 5253 29687 5287
rect 29687 5253 29696 5287
rect 29644 5244 29696 5253
rect 29736 5287 29788 5296
rect 29736 5253 29745 5287
rect 29745 5253 29779 5287
rect 29779 5253 29788 5287
rect 29736 5244 29788 5253
rect 26516 5219 26568 5228
rect 26516 5185 26525 5219
rect 26525 5185 26559 5219
rect 26559 5185 26568 5219
rect 26516 5176 26568 5185
rect 18236 5108 18288 5160
rect 21640 5108 21692 5160
rect 22560 5151 22612 5160
rect 22560 5117 22569 5151
rect 22569 5117 22603 5151
rect 22603 5117 22612 5151
rect 22560 5108 22612 5117
rect 23204 5151 23256 5160
rect 23204 5117 23213 5151
rect 23213 5117 23247 5151
rect 23247 5117 23256 5151
rect 23204 5108 23256 5117
rect 24860 5151 24912 5160
rect 24860 5117 24869 5151
rect 24869 5117 24903 5151
rect 24903 5117 24912 5151
rect 24860 5108 24912 5117
rect 27252 5151 27304 5160
rect 27252 5117 27261 5151
rect 27261 5117 27295 5151
rect 27295 5117 27304 5151
rect 27252 5108 27304 5117
rect 27620 5151 27672 5160
rect 27620 5117 27629 5151
rect 27629 5117 27663 5151
rect 27663 5117 27672 5151
rect 27620 5108 27672 5117
rect 28816 5151 28868 5160
rect 28816 5117 28825 5151
rect 28825 5117 28859 5151
rect 28859 5117 28868 5151
rect 28816 5108 28868 5117
rect 21180 4972 21232 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 18236 4811 18288 4820
rect 18236 4777 18245 4811
rect 18245 4777 18279 4811
rect 18279 4777 18288 4811
rect 18236 4768 18288 4777
rect 22560 4768 22612 4820
rect 27252 4768 27304 4820
rect 28264 4768 28316 4820
rect 21180 4675 21232 4684
rect 21180 4641 21189 4675
rect 21189 4641 21223 4675
rect 21223 4641 21232 4675
rect 21180 4632 21232 4641
rect 21824 4675 21876 4684
rect 21824 4641 21833 4675
rect 21833 4641 21867 4675
rect 21867 4641 21876 4675
rect 21824 4632 21876 4641
rect 19340 4564 19392 4616
rect 20352 4607 20404 4616
rect 20352 4573 20361 4607
rect 20361 4573 20395 4607
rect 20395 4573 20404 4607
rect 20352 4564 20404 4573
rect 22836 4607 22888 4616
rect 22836 4573 22845 4607
rect 22845 4573 22879 4607
rect 22879 4573 22888 4607
rect 22836 4564 22888 4573
rect 25504 4632 25556 4684
rect 25964 4675 26016 4684
rect 25964 4641 25973 4675
rect 25973 4641 26007 4675
rect 26007 4641 26016 4675
rect 25964 4632 26016 4641
rect 29000 4632 29052 4684
rect 29276 4564 29328 4616
rect 30104 4564 30156 4616
rect 20352 4428 20404 4480
rect 23480 4496 23532 4548
rect 25044 4496 25096 4548
rect 25412 4539 25464 4548
rect 25412 4505 25421 4539
rect 25421 4505 25455 4539
rect 25455 4505 25464 4539
rect 25412 4496 25464 4505
rect 26424 4428 26476 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 20352 4131 20404 4140
rect 20352 4097 20361 4131
rect 20361 4097 20395 4131
rect 20395 4097 20404 4131
rect 20352 4088 20404 4097
rect 22836 4224 22888 4276
rect 25412 4267 25464 4276
rect 25412 4233 25421 4267
rect 25421 4233 25455 4267
rect 25455 4233 25464 4267
rect 25412 4224 25464 4233
rect 21456 4088 21508 4140
rect 23480 4156 23532 4208
rect 25504 4131 25556 4140
rect 25504 4097 25513 4131
rect 25513 4097 25547 4131
rect 25547 4097 25556 4131
rect 25504 4088 25556 4097
rect 26516 4131 26568 4140
rect 26516 4097 26525 4131
rect 26525 4097 26559 4131
rect 26559 4097 26568 4131
rect 26516 4088 26568 4097
rect 29184 4088 29236 4140
rect 22284 4020 22336 4072
rect 24124 4063 24176 4072
rect 18604 3952 18656 4004
rect 24124 4029 24133 4063
rect 24133 4029 24167 4063
rect 24167 4029 24176 4063
rect 24124 4020 24176 4029
rect 26884 4020 26936 4072
rect 16120 3927 16172 3936
rect 16120 3893 16129 3927
rect 16129 3893 16163 3927
rect 16163 3893 16172 3927
rect 16120 3884 16172 3893
rect 17224 3927 17276 3936
rect 17224 3893 17233 3927
rect 17233 3893 17267 3927
rect 17267 3893 17276 3927
rect 17224 3884 17276 3893
rect 19432 3884 19484 3936
rect 21272 3884 21324 3936
rect 23756 3884 23808 3936
rect 28724 3884 28776 3936
rect 30196 3927 30248 3936
rect 30196 3893 30205 3927
rect 30205 3893 30239 3927
rect 30239 3893 30248 3927
rect 30196 3884 30248 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 20076 3680 20128 3732
rect 16856 3612 16908 3664
rect 19156 3612 19208 3664
rect 19340 3612 19392 3664
rect 31024 3612 31076 3664
rect 17776 3544 17828 3596
rect 22744 3587 22796 3596
rect 22744 3553 22753 3587
rect 22753 3553 22787 3587
rect 22787 3553 22796 3587
rect 22744 3544 22796 3553
rect 28540 3587 28592 3596
rect 28540 3553 28549 3587
rect 28549 3553 28583 3587
rect 28583 3553 28592 3587
rect 28540 3544 28592 3553
rect 30196 3544 30248 3596
rect 4160 3476 4212 3528
rect 5172 3519 5224 3528
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 5172 3476 5224 3485
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 6828 3519 6880 3528
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 11796 3476 11848 3528
rect 12532 3476 12584 3528
rect 13084 3476 13136 3528
rect 13636 3519 13688 3528
rect 13636 3485 13645 3519
rect 13645 3485 13679 3519
rect 13679 3485 13688 3519
rect 13636 3476 13688 3485
rect 15016 3519 15068 3528
rect 15016 3485 15025 3519
rect 15025 3485 15059 3519
rect 15059 3485 15068 3519
rect 15016 3476 15068 3485
rect 16396 3476 16448 3528
rect 21548 3519 21600 3528
rect 21548 3485 21557 3519
rect 21557 3485 21591 3519
rect 21591 3485 21600 3519
rect 21548 3476 21600 3485
rect 25504 3476 25556 3528
rect 26516 3519 26568 3528
rect 26516 3485 26525 3519
rect 26525 3485 26559 3519
rect 26559 3485 26568 3519
rect 26516 3476 26568 3485
rect 29736 3519 29788 3528
rect 29736 3485 29745 3519
rect 29745 3485 29779 3519
rect 29779 3485 29788 3519
rect 29736 3476 29788 3485
rect 29920 3476 29972 3528
rect 30472 3476 30524 3528
rect 31852 3476 31904 3528
rect 32680 3476 32732 3528
rect 33232 3476 33284 3528
rect 35348 3476 35400 3528
rect 35440 3476 35492 3528
rect 36268 3519 36320 3528
rect 36268 3485 36277 3519
rect 36277 3485 36311 3519
rect 36311 3485 36320 3519
rect 36268 3476 36320 3485
rect 37096 3519 37148 3528
rect 37096 3485 37105 3519
rect 37105 3485 37139 3519
rect 37139 3485 37148 3519
rect 37096 3476 37148 3485
rect 37924 3519 37976 3528
rect 37924 3485 37933 3519
rect 37933 3485 37967 3519
rect 37967 3485 37976 3519
rect 37924 3476 37976 3485
rect 39028 3519 39080 3528
rect 39028 3485 39037 3519
rect 39037 3485 39071 3519
rect 39071 3485 39080 3519
rect 39028 3476 39080 3485
rect 40408 3519 40460 3528
rect 40408 3485 40417 3519
rect 40417 3485 40451 3519
rect 40451 3485 40460 3519
rect 40408 3476 40460 3485
rect 40960 3476 41012 3528
rect 41512 3519 41564 3528
rect 41512 3485 41521 3519
rect 41521 3485 41555 3519
rect 41555 3485 41564 3519
rect 41512 3476 41564 3485
rect 42892 3519 42944 3528
rect 42892 3485 42901 3519
rect 42901 3485 42935 3519
rect 42935 3485 42944 3519
rect 42892 3476 42944 3485
rect 43168 3476 43220 3528
rect 44824 3476 44876 3528
rect 45652 3476 45704 3528
rect 46480 3519 46532 3528
rect 46480 3485 46489 3519
rect 46489 3485 46523 3519
rect 46523 3485 46532 3519
rect 46480 3476 46532 3485
rect 46756 3476 46808 3528
rect 47308 3476 47360 3528
rect 18880 3408 18932 3460
rect 20168 3451 20220 3460
rect 20168 3417 20177 3451
rect 20177 3417 20211 3451
rect 20211 3417 20220 3451
rect 20168 3408 20220 3417
rect 21364 3408 21416 3460
rect 28724 3451 28776 3460
rect 28724 3417 28733 3451
rect 28733 3417 28767 3451
rect 28767 3417 28776 3451
rect 28724 3408 28776 3417
rect 29644 3408 29696 3460
rect 30840 3408 30892 3460
rect 25412 3383 25464 3392
rect 25412 3349 25421 3383
rect 25421 3349 25455 3383
rect 25455 3349 25464 3383
rect 25412 3340 25464 3349
rect 28080 3340 28132 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 20168 3136 20220 3188
rect 20536 3068 20588 3120
rect 22192 3111 22244 3120
rect 22192 3077 22201 3111
rect 22201 3077 22235 3111
rect 22235 3077 22244 3111
rect 22192 3068 22244 3077
rect 23756 3068 23808 3120
rect 25412 3111 25464 3120
rect 25412 3077 25421 3111
rect 25421 3077 25455 3111
rect 25455 3077 25464 3111
rect 25412 3068 25464 3077
rect 28080 3111 28132 3120
rect 28080 3077 28089 3111
rect 28089 3077 28123 3111
rect 28123 3077 28132 3111
rect 28080 3068 28132 3077
rect 18880 3043 18932 3052
rect 18880 3009 18889 3043
rect 18889 3009 18923 3043
rect 18923 3009 18932 3043
rect 18880 3000 18932 3009
rect 20352 3043 20404 3052
rect 20352 3009 20361 3043
rect 20361 3009 20395 3043
rect 20395 3009 20404 3043
rect 20352 3000 20404 3009
rect 21548 3000 21600 3052
rect 30104 3000 30156 3052
rect 5448 2932 5500 2984
rect 7932 2932 7984 2984
rect 9864 2932 9916 2984
rect 15292 2932 15344 2984
rect 17500 2932 17552 2984
rect 4896 2864 4948 2916
rect 6276 2864 6328 2916
rect 3148 2796 3200 2848
rect 3884 2796 3936 2848
rect 6552 2796 6604 2848
rect 8760 2864 8812 2916
rect 11244 2864 11296 2916
rect 13360 2864 13412 2916
rect 14464 2864 14516 2916
rect 18052 2864 18104 2916
rect 9036 2796 9088 2848
rect 10692 2796 10744 2848
rect 12072 2796 12124 2848
rect 13912 2796 13964 2848
rect 15844 2796 15896 2848
rect 19340 2932 19392 2984
rect 22468 2975 22520 2984
rect 22468 2941 22477 2975
rect 22477 2941 22511 2975
rect 22511 2941 22520 2975
rect 22468 2932 22520 2941
rect 24400 2975 24452 2984
rect 24400 2941 24409 2975
rect 24409 2941 24443 2975
rect 24443 2941 24452 2975
rect 24400 2932 24452 2941
rect 24584 2932 24636 2984
rect 25780 2975 25832 2984
rect 25780 2941 25789 2975
rect 25789 2941 25823 2975
rect 25823 2941 25832 2975
rect 25780 2932 25832 2941
rect 27160 2975 27212 2984
rect 27160 2941 27169 2975
rect 27169 2941 27203 2975
rect 27203 2941 27212 2975
rect 27160 2932 27212 2941
rect 29184 2932 29236 2984
rect 29368 2975 29420 2984
rect 29368 2941 29377 2975
rect 29377 2941 29411 2975
rect 29411 2941 29420 2975
rect 29368 2932 29420 2941
rect 31208 2932 31260 2984
rect 32956 2932 33008 2984
rect 38752 2932 38804 2984
rect 40684 2932 40736 2984
rect 42616 2932 42668 2984
rect 44548 2932 44600 2984
rect 34796 2864 34848 2916
rect 19984 2796 20036 2848
rect 22836 2796 22888 2848
rect 30196 2796 30248 2848
rect 31300 2796 31352 2848
rect 32404 2796 32456 2848
rect 33784 2796 33836 2848
rect 34336 2796 34388 2848
rect 35716 2796 35768 2848
rect 36820 2796 36872 2848
rect 37648 2796 37700 2848
rect 38200 2796 38252 2848
rect 39580 2796 39632 2848
rect 40132 2796 40184 2848
rect 42064 2796 42116 2848
rect 43444 2796 43496 2848
rect 43996 2796 44048 2848
rect 45376 2796 45428 2848
rect 45928 2796 45980 2848
rect 47032 2796 47084 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 19340 2592 19392 2644
rect 22192 2592 22244 2644
rect 26424 2635 26476 2644
rect 26424 2601 26433 2635
rect 26433 2601 26467 2635
rect 26467 2601 26476 2635
rect 26424 2592 26476 2601
rect 29184 2592 29236 2644
rect 31208 2635 31260 2644
rect 31208 2601 31217 2635
rect 31217 2601 31251 2635
rect 31251 2601 31260 2635
rect 31208 2592 31260 2601
rect 7104 2524 7156 2576
rect 9588 2524 9640 2576
rect 11520 2524 11572 2576
rect 14188 2524 14240 2576
rect 20260 2524 20312 2576
rect 3516 2456 3568 2508
rect 8208 2456 8260 2508
rect 10416 2456 10468 2508
rect 12808 2456 12860 2508
rect 14740 2456 14792 2508
rect 16672 2456 16724 2508
rect 2596 2388 2648 2440
rect 4620 2388 4672 2440
rect 5724 2388 5776 2440
rect 12256 2388 12308 2440
rect 15568 2388 15620 2440
rect 18880 2456 18932 2508
rect 23020 2499 23072 2508
rect 23020 2465 23029 2499
rect 23029 2465 23063 2499
rect 23063 2465 23072 2499
rect 23020 2456 23072 2465
rect 32128 2524 32180 2576
rect 34612 2524 34664 2576
rect 38476 2524 38528 2576
rect 42340 2524 42392 2576
rect 45100 2524 45152 2576
rect 25504 2499 25556 2508
rect 25504 2465 25513 2499
rect 25513 2465 25547 2499
rect 25547 2465 25556 2499
rect 25504 2456 25556 2465
rect 28264 2499 28316 2508
rect 28264 2465 28273 2499
rect 28273 2465 28307 2499
rect 28307 2465 28316 2499
rect 28264 2456 28316 2465
rect 29736 2456 29788 2508
rect 31576 2456 31628 2508
rect 33508 2456 33560 2508
rect 36544 2456 36596 2508
rect 39304 2456 39356 2508
rect 41236 2456 41288 2508
rect 43720 2456 43772 2508
rect 7380 2320 7432 2372
rect 20812 2388 20864 2440
rect 30104 2431 30156 2440
rect 18328 2320 18380 2372
rect 20352 2320 20404 2372
rect 30104 2397 30113 2431
rect 30113 2397 30147 2431
rect 30147 2397 30156 2431
rect 30104 2388 30156 2397
rect 30748 2388 30800 2440
rect 34060 2388 34112 2440
rect 35992 2388 36044 2440
rect 22836 2363 22888 2372
rect 22836 2329 22845 2363
rect 22845 2329 22879 2363
rect 22879 2329 22888 2363
rect 25044 2363 25096 2372
rect 22836 2320 22888 2329
rect 25044 2329 25053 2363
rect 25053 2329 25087 2363
rect 25087 2329 25096 2363
rect 25044 2320 25096 2329
rect 24584 2252 24636 2304
rect 37372 2320 37424 2372
rect 39856 2388 39908 2440
rect 41788 2388 41840 2440
rect 44272 2320 44324 2372
rect 46204 2388 46256 2440
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 3974 49200 4030 50000
rect 4342 49200 4398 50000
rect 4710 49200 4766 50000
rect 5078 49314 5134 50000
rect 4816 49286 5134 49314
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4724 47258 4752 49200
rect 4712 47252 4764 47258
rect 4712 47194 4764 47200
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4816 45554 4844 49286
rect 5078 49200 5134 49286
rect 5446 49200 5502 50000
rect 5814 49200 5870 50000
rect 6182 49314 6238 50000
rect 6012 49286 6238 49314
rect 5828 47258 5856 49200
rect 6012 47258 6040 49286
rect 6182 49200 6238 49286
rect 6550 49200 6606 50000
rect 6918 49200 6974 50000
rect 7286 49314 7342 50000
rect 7116 49286 7342 49314
rect 5816 47252 5868 47258
rect 5816 47194 5868 47200
rect 6000 47252 6052 47258
rect 6000 47194 6052 47200
rect 6932 46578 6960 49200
rect 7116 47258 7144 49286
rect 7286 49200 7342 49286
rect 7654 49200 7710 50000
rect 8022 49314 8078 50000
rect 7760 49286 8078 49314
rect 7760 47258 7788 49286
rect 8022 49200 8078 49286
rect 8390 49200 8446 50000
rect 8758 49200 8814 50000
rect 9126 49200 9182 50000
rect 9494 49200 9550 50000
rect 9862 49200 9918 50000
rect 10230 49200 10286 50000
rect 10598 49200 10654 50000
rect 10966 49200 11022 50000
rect 11334 49314 11390 50000
rect 11164 49286 11390 49314
rect 8404 47258 8432 49200
rect 9140 47258 9168 49200
rect 7104 47252 7156 47258
rect 7104 47194 7156 47200
rect 7748 47252 7800 47258
rect 7748 47194 7800 47200
rect 8392 47252 8444 47258
rect 8392 47194 8444 47200
rect 9128 47252 9180 47258
rect 9128 47194 9180 47200
rect 9508 46646 9536 49200
rect 10244 47258 10272 49200
rect 10232 47252 10284 47258
rect 10232 47194 10284 47200
rect 10612 46918 10640 49200
rect 11164 47258 11192 49286
rect 11334 49200 11390 49286
rect 11702 49200 11758 50000
rect 12070 49200 12126 50000
rect 12438 49200 12494 50000
rect 12806 49200 12862 50000
rect 13174 49200 13230 50000
rect 13542 49200 13598 50000
rect 13910 49200 13966 50000
rect 14278 49200 14334 50000
rect 14646 49200 14702 50000
rect 15014 49200 15070 50000
rect 15382 49200 15438 50000
rect 15750 49314 15806 50000
rect 15580 49286 15806 49314
rect 11152 47252 11204 47258
rect 11152 47194 11204 47200
rect 10600 46912 10652 46918
rect 10600 46854 10652 46860
rect 9496 46640 9548 46646
rect 9496 46582 9548 46588
rect 6920 46572 6972 46578
rect 6920 46514 6972 46520
rect 11716 46170 11744 49200
rect 12452 47258 12480 49200
rect 12440 47252 12492 47258
rect 12440 47194 12492 47200
rect 11704 46164 11756 46170
rect 11704 46106 11756 46112
rect 12820 45898 12848 49200
rect 13556 47258 13584 49200
rect 13544 47252 13596 47258
rect 13544 47194 13596 47200
rect 13924 46510 13952 49200
rect 14660 46578 14688 49200
rect 14648 46572 14700 46578
rect 14648 46514 14700 46520
rect 13912 46504 13964 46510
rect 13912 46446 13964 46452
rect 15028 46442 15056 49200
rect 15580 46578 15608 49286
rect 15750 49200 15806 49286
rect 16118 49200 16174 50000
rect 16486 49200 16542 50000
rect 16854 49200 16910 50000
rect 17222 49200 17278 50000
rect 17590 49200 17646 50000
rect 17958 49200 18014 50000
rect 18326 49314 18382 50000
rect 18326 49286 18644 49314
rect 18326 49200 18382 49286
rect 16132 46714 16160 49200
rect 16868 47258 16896 49200
rect 16856 47252 16908 47258
rect 16856 47194 16908 47200
rect 17132 46912 17184 46918
rect 17132 46854 17184 46860
rect 16120 46708 16172 46714
rect 16120 46650 16172 46656
rect 15568 46572 15620 46578
rect 15568 46514 15620 46520
rect 15016 46436 15068 46442
rect 15016 46378 15068 46384
rect 16132 46102 16160 46650
rect 16120 46096 16172 46102
rect 16120 46038 16172 46044
rect 12808 45892 12860 45898
rect 12808 45834 12860 45840
rect 17144 45626 17172 46854
rect 17236 46714 17264 49200
rect 17224 46708 17276 46714
rect 17224 46650 17276 46656
rect 17408 46572 17460 46578
rect 17408 46514 17460 46520
rect 17420 45966 17448 46514
rect 17592 46504 17644 46510
rect 17592 46446 17644 46452
rect 17604 46170 17632 46446
rect 17592 46164 17644 46170
rect 17592 46106 17644 46112
rect 17408 45960 17460 45966
rect 17408 45902 17460 45908
rect 17132 45620 17184 45626
rect 17132 45562 17184 45568
rect 4632 45526 4844 45554
rect 4632 45422 4660 45526
rect 17972 45490 18000 49200
rect 18144 46980 18196 46986
rect 18144 46922 18196 46928
rect 18052 46572 18104 46578
rect 18052 46514 18104 46520
rect 17960 45484 18012 45490
rect 17960 45426 18012 45432
rect 4620 45416 4672 45422
rect 4620 45358 4672 45364
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 18064 44470 18092 46514
rect 18156 44878 18184 46922
rect 18616 46918 18644 49286
rect 18694 49200 18750 50000
rect 19062 49200 19118 50000
rect 19430 49200 19486 50000
rect 19798 49200 19854 50000
rect 20166 49200 20222 50000
rect 20534 49200 20590 50000
rect 20902 49200 20958 50000
rect 21270 49200 21326 50000
rect 21638 49200 21694 50000
rect 22006 49200 22062 50000
rect 22374 49200 22430 50000
rect 22742 49200 22798 50000
rect 23110 49200 23166 50000
rect 23478 49450 23534 50000
rect 23478 49422 23704 49450
rect 23478 49200 23534 49422
rect 18696 47048 18748 47054
rect 18696 46990 18748 46996
rect 18420 46912 18472 46918
rect 18420 46854 18472 46860
rect 18604 46912 18656 46918
rect 18604 46854 18656 46860
rect 18432 46578 18460 46854
rect 18328 46572 18380 46578
rect 18328 46514 18380 46520
rect 18420 46572 18472 46578
rect 18420 46514 18472 46520
rect 18340 45082 18368 46514
rect 18604 46504 18656 46510
rect 18708 46458 18736 46990
rect 18972 46980 19024 46986
rect 18972 46922 19024 46928
rect 18984 46617 19012 46922
rect 18970 46608 19026 46617
rect 18970 46543 18972 46552
rect 19024 46543 19026 46552
rect 18972 46514 19024 46520
rect 18656 46452 18736 46458
rect 18604 46446 18736 46452
rect 18616 46430 18736 46446
rect 18708 46170 18736 46430
rect 18788 46368 18840 46374
rect 18788 46310 18840 46316
rect 18696 46164 18748 46170
rect 18696 46106 18748 46112
rect 18800 45490 18828 46310
rect 18788 45484 18840 45490
rect 18788 45426 18840 45432
rect 18972 45484 19024 45490
rect 18972 45426 19024 45432
rect 18328 45076 18380 45082
rect 18328 45018 18380 45024
rect 18144 44872 18196 44878
rect 18144 44814 18196 44820
rect 18800 44742 18828 45426
rect 18788 44736 18840 44742
rect 18788 44678 18840 44684
rect 18984 44538 19012 45426
rect 18972 44532 19024 44538
rect 18972 44474 19024 44480
rect 18052 44464 18104 44470
rect 18052 44406 18104 44412
rect 19076 44402 19104 49200
rect 19444 46510 19472 49200
rect 19708 47796 19760 47802
rect 19708 47738 19760 47744
rect 19720 47190 19748 47738
rect 20180 47258 20208 49200
rect 20168 47252 20220 47258
rect 20168 47194 20220 47200
rect 19708 47184 19760 47190
rect 19708 47126 19760 47132
rect 19892 47184 19944 47190
rect 19892 47126 19944 47132
rect 19904 47054 19932 47126
rect 19892 47048 19944 47054
rect 20444 47048 20496 47054
rect 19944 47008 20024 47036
rect 19892 46990 19944 46996
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19996 46646 20024 47008
rect 20444 46990 20496 46996
rect 19984 46640 20036 46646
rect 19984 46582 20036 46588
rect 20456 46578 20484 46990
rect 19892 46572 19944 46578
rect 19892 46514 19944 46520
rect 20444 46572 20496 46578
rect 20444 46514 20496 46520
rect 19432 46504 19484 46510
rect 19338 46472 19394 46481
rect 19904 46458 19932 46514
rect 19432 46446 19484 46452
rect 19338 46407 19340 46416
rect 19392 46407 19394 46416
rect 19812 46430 19932 46458
rect 19340 46378 19392 46384
rect 19432 46368 19484 46374
rect 19432 46310 19484 46316
rect 19340 46028 19392 46034
rect 19340 45970 19392 45976
rect 19352 45626 19380 45970
rect 19444 45830 19472 46310
rect 19812 45966 19840 46430
rect 19984 46368 20036 46374
rect 19984 46310 20036 46316
rect 19800 45960 19852 45966
rect 19800 45902 19852 45908
rect 19892 45960 19944 45966
rect 19892 45902 19944 45908
rect 19904 45830 19932 45902
rect 19432 45824 19484 45830
rect 19432 45766 19484 45772
rect 19892 45824 19944 45830
rect 19892 45766 19944 45772
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19340 45620 19392 45626
rect 19340 45562 19392 45568
rect 19996 44878 20024 46310
rect 20548 45626 20576 49200
rect 20628 47252 20680 47258
rect 20628 47194 20680 47200
rect 20640 45830 20668 47194
rect 21180 46912 21232 46918
rect 21180 46854 21232 46860
rect 20904 46504 20956 46510
rect 20904 46446 20956 46452
rect 20916 46345 20944 46446
rect 20902 46336 20958 46345
rect 20902 46271 20958 46280
rect 21192 46102 21220 46854
rect 21180 46096 21232 46102
rect 21180 46038 21232 46044
rect 21088 45892 21140 45898
rect 21088 45834 21140 45840
rect 20628 45824 20680 45830
rect 20628 45766 20680 45772
rect 20640 45626 20668 45766
rect 20536 45620 20588 45626
rect 20536 45562 20588 45568
rect 20628 45620 20680 45626
rect 20628 45562 20680 45568
rect 20168 45416 20220 45422
rect 20168 45358 20220 45364
rect 19984 44872 20036 44878
rect 19984 44814 20036 44820
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19996 44402 20024 44814
rect 19064 44396 19116 44402
rect 19064 44338 19116 44344
rect 19984 44396 20036 44402
rect 19984 44338 20036 44344
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 20180 43858 20208 45358
rect 20548 44538 20576 45562
rect 20640 45354 20668 45562
rect 20904 45484 20956 45490
rect 20904 45426 20956 45432
rect 20996 45484 21048 45490
rect 20996 45426 21048 45432
rect 20628 45348 20680 45354
rect 20628 45290 20680 45296
rect 20536 44532 20588 44538
rect 20536 44474 20588 44480
rect 20536 44396 20588 44402
rect 20536 44338 20588 44344
rect 20548 43926 20576 44338
rect 20536 43920 20588 43926
rect 20536 43862 20588 43868
rect 20168 43852 20220 43858
rect 20168 43794 20220 43800
rect 20548 43790 20576 43862
rect 20536 43784 20588 43790
rect 20536 43726 20588 43732
rect 20640 43654 20668 45290
rect 20916 44946 20944 45426
rect 20904 44940 20956 44946
rect 20904 44882 20956 44888
rect 21008 44878 21036 45426
rect 20996 44872 21048 44878
rect 20996 44814 21048 44820
rect 21100 44402 21128 45834
rect 21088 44396 21140 44402
rect 21088 44338 21140 44344
rect 20720 44328 20772 44334
rect 20720 44270 20772 44276
rect 20732 43790 20760 44270
rect 20720 43784 20772 43790
rect 20720 43726 20772 43732
rect 20628 43648 20680 43654
rect 20628 43590 20680 43596
rect 21180 43648 21232 43654
rect 21180 43590 21232 43596
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 21192 41414 21220 43590
rect 21284 43314 21312 49200
rect 21456 46912 21508 46918
rect 21456 46854 21508 46860
rect 21468 46510 21496 46854
rect 21652 46714 21680 49200
rect 22388 47802 22416 49200
rect 22376 47796 22428 47802
rect 22376 47738 22428 47744
rect 22100 47048 22152 47054
rect 22100 46990 22152 46996
rect 22112 46753 22140 46990
rect 21822 46744 21878 46753
rect 21640 46708 21692 46714
rect 21822 46679 21878 46688
rect 22098 46744 22154 46753
rect 22098 46679 22154 46688
rect 21640 46650 21692 46656
rect 21732 46640 21784 46646
rect 21732 46582 21784 46588
rect 21456 46504 21508 46510
rect 21456 46446 21508 46452
rect 21744 45966 21772 46582
rect 21836 45966 21864 46679
rect 22100 46572 22152 46578
rect 22100 46514 22152 46520
rect 22112 46345 22140 46514
rect 22756 46442 22784 49200
rect 22836 46572 22888 46578
rect 22836 46514 22888 46520
rect 22848 46481 22876 46514
rect 22834 46472 22890 46481
rect 22744 46436 22796 46442
rect 22834 46407 22890 46416
rect 22744 46378 22796 46384
rect 22098 46336 22154 46345
rect 22098 46271 22154 46280
rect 22756 45966 22784 46378
rect 21732 45960 21784 45966
rect 21732 45902 21784 45908
rect 21824 45960 21876 45966
rect 21824 45902 21876 45908
rect 22744 45960 22796 45966
rect 22744 45902 22796 45908
rect 23204 45960 23256 45966
rect 23204 45902 23256 45908
rect 21744 43994 21772 45902
rect 23112 45892 23164 45898
rect 23112 45834 23164 45840
rect 23124 45422 23152 45834
rect 23216 45490 23244 45902
rect 23480 45552 23532 45558
rect 23480 45494 23532 45500
rect 23204 45484 23256 45490
rect 23204 45426 23256 45432
rect 23020 45416 23072 45422
rect 23020 45358 23072 45364
rect 23112 45416 23164 45422
rect 23112 45358 23164 45364
rect 23032 44878 23060 45358
rect 23124 45014 23152 45358
rect 23112 45008 23164 45014
rect 23112 44950 23164 44956
rect 22008 44872 22060 44878
rect 22008 44814 22060 44820
rect 23020 44872 23072 44878
rect 23020 44814 23072 44820
rect 21916 44736 21968 44742
rect 21916 44678 21968 44684
rect 21928 44470 21956 44678
rect 22020 44538 22048 44814
rect 22192 44804 22244 44810
rect 22192 44746 22244 44752
rect 22008 44532 22060 44538
rect 22008 44474 22060 44480
rect 21916 44464 21968 44470
rect 21916 44406 21968 44412
rect 21732 43988 21784 43994
rect 21732 43930 21784 43936
rect 21928 43858 21956 44406
rect 21916 43852 21968 43858
rect 21916 43794 21968 43800
rect 21272 43308 21324 43314
rect 21272 43250 21324 43256
rect 22020 43246 22048 44474
rect 22204 43314 22232 44746
rect 22376 44736 22428 44742
rect 22376 44678 22428 44684
rect 22388 44538 22416 44678
rect 22376 44532 22428 44538
rect 22376 44474 22428 44480
rect 23032 44470 23060 44814
rect 23124 44538 23152 44950
rect 23112 44532 23164 44538
rect 23112 44474 23164 44480
rect 22652 44464 22704 44470
rect 22836 44464 22888 44470
rect 22704 44424 22836 44452
rect 22652 44406 22704 44412
rect 22836 44406 22888 44412
rect 23020 44464 23072 44470
rect 23020 44406 23072 44412
rect 22928 44396 22980 44402
rect 22928 44338 22980 44344
rect 22744 43784 22796 43790
rect 22940 43772 22968 44338
rect 23112 44328 23164 44334
rect 23112 44270 23164 44276
rect 22796 43744 22968 43772
rect 22744 43726 22796 43732
rect 22192 43308 22244 43314
rect 22192 43250 22244 43256
rect 22008 43240 22060 43246
rect 22008 43182 22060 43188
rect 22020 42022 22048 43182
rect 22652 42696 22704 42702
rect 22652 42638 22704 42644
rect 22664 42362 22692 42638
rect 22940 42566 22968 43744
rect 23124 43722 23152 44270
rect 23112 43716 23164 43722
rect 23112 43658 23164 43664
rect 23020 43648 23072 43654
rect 23020 43590 23072 43596
rect 23032 42702 23060 43590
rect 23124 43382 23152 43658
rect 23112 43376 23164 43382
rect 23112 43318 23164 43324
rect 23216 42906 23244 45426
rect 23492 44878 23520 45494
rect 23480 44872 23532 44878
rect 23480 44814 23532 44820
rect 23296 43716 23348 43722
rect 23296 43658 23348 43664
rect 23388 43716 23440 43722
rect 23388 43658 23440 43664
rect 23308 43246 23336 43658
rect 23400 43314 23428 43658
rect 23388 43308 23440 43314
rect 23388 43250 23440 43256
rect 23296 43240 23348 43246
rect 23296 43182 23348 43188
rect 23676 43178 23704 49422
rect 23846 49200 23902 50000
rect 24214 49200 24270 50000
rect 24582 49314 24638 50000
rect 24412 49286 24638 49314
rect 23860 46646 23888 49200
rect 24228 46918 24256 49200
rect 24216 46912 24268 46918
rect 24216 46854 24268 46860
rect 23848 46640 23900 46646
rect 23848 46582 23900 46588
rect 23860 45626 23888 46582
rect 24124 46572 24176 46578
rect 24124 46514 24176 46520
rect 24308 46572 24360 46578
rect 24308 46514 24360 46520
rect 23848 45620 23900 45626
rect 23848 45562 23900 45568
rect 24136 44946 24164 46514
rect 24320 46034 24348 46514
rect 24308 46028 24360 46034
rect 24308 45970 24360 45976
rect 24308 45620 24360 45626
rect 24308 45562 24360 45568
rect 24216 45280 24268 45286
rect 24216 45222 24268 45228
rect 24124 44940 24176 44946
rect 24124 44882 24176 44888
rect 24228 44878 24256 45222
rect 24216 44872 24268 44878
rect 24216 44814 24268 44820
rect 24228 44538 24256 44814
rect 24320 44742 24348 45562
rect 24308 44736 24360 44742
rect 24308 44678 24360 44684
rect 24216 44532 24268 44538
rect 24216 44474 24268 44480
rect 24320 44402 24348 44678
rect 24308 44396 24360 44402
rect 24308 44338 24360 44344
rect 24412 43994 24440 49286
rect 24582 49200 24638 49286
rect 24950 49200 25006 50000
rect 25318 49200 25374 50000
rect 25686 49200 25742 50000
rect 26054 49200 26110 50000
rect 26422 49314 26478 50000
rect 26422 49286 26648 49314
rect 26422 49200 26478 49286
rect 24860 46368 24912 46374
rect 24860 46310 24912 46316
rect 24872 46170 24900 46310
rect 24860 46164 24912 46170
rect 24860 46106 24912 46112
rect 24768 46096 24820 46102
rect 24768 46038 24820 46044
rect 24584 45892 24636 45898
rect 24584 45834 24636 45840
rect 24596 45558 24624 45834
rect 24584 45552 24636 45558
rect 24584 45494 24636 45500
rect 24780 44402 24808 46038
rect 24964 45082 24992 49200
rect 25136 47048 25188 47054
rect 25136 46990 25188 46996
rect 25148 45558 25176 46990
rect 25332 45558 25360 49200
rect 25700 47258 25728 49200
rect 26068 47258 26096 49200
rect 25688 47252 25740 47258
rect 25688 47194 25740 47200
rect 26056 47252 26108 47258
rect 26056 47194 26108 47200
rect 25596 47048 25648 47054
rect 25596 46990 25648 46996
rect 25608 46578 25636 46990
rect 26424 46912 26476 46918
rect 26424 46854 26476 46860
rect 25596 46572 25648 46578
rect 25596 46514 25648 46520
rect 25412 46436 25464 46442
rect 25412 46378 25464 46384
rect 25424 45830 25452 46378
rect 25412 45824 25464 45830
rect 25412 45766 25464 45772
rect 25136 45552 25188 45558
rect 25136 45494 25188 45500
rect 25320 45552 25372 45558
rect 25320 45494 25372 45500
rect 25228 45280 25280 45286
rect 25228 45222 25280 45228
rect 24952 45076 25004 45082
rect 24952 45018 25004 45024
rect 25240 44402 25268 45222
rect 25332 44878 25360 45494
rect 25412 45484 25464 45490
rect 25412 45426 25464 45432
rect 25424 44946 25452 45426
rect 25504 45348 25556 45354
rect 25504 45290 25556 45296
rect 25516 45082 25544 45290
rect 25504 45076 25556 45082
rect 25504 45018 25556 45024
rect 25608 45014 25636 46514
rect 26436 46510 26464 46854
rect 26424 46504 26476 46510
rect 26424 46446 26476 46452
rect 26240 46368 26292 46374
rect 26240 46310 26292 46316
rect 26148 46028 26200 46034
rect 26148 45970 26200 45976
rect 26056 45960 26108 45966
rect 26056 45902 26108 45908
rect 26068 45490 26096 45902
rect 26160 45490 26188 45970
rect 26252 45966 26280 46310
rect 26240 45960 26292 45966
rect 26240 45902 26292 45908
rect 26332 45960 26384 45966
rect 26332 45902 26384 45908
rect 26056 45484 26108 45490
rect 26056 45426 26108 45432
rect 26148 45484 26200 45490
rect 26148 45426 26200 45432
rect 26068 45014 26096 45426
rect 25596 45008 25648 45014
rect 25596 44950 25648 44956
rect 26056 45008 26108 45014
rect 26056 44950 26108 44956
rect 25412 44940 25464 44946
rect 25412 44882 25464 44888
rect 25320 44872 25372 44878
rect 25320 44814 25372 44820
rect 25964 44872 26016 44878
rect 25964 44814 26016 44820
rect 24768 44396 24820 44402
rect 24768 44338 24820 44344
rect 25228 44396 25280 44402
rect 25228 44338 25280 44344
rect 24400 43988 24452 43994
rect 24400 43930 24452 43936
rect 24780 43790 24808 44338
rect 24768 43784 24820 43790
rect 24768 43726 24820 43732
rect 24584 43376 24636 43382
rect 24584 43318 24636 43324
rect 23756 43308 23808 43314
rect 23756 43250 23808 43256
rect 24032 43308 24084 43314
rect 24032 43250 24084 43256
rect 23664 43172 23716 43178
rect 23664 43114 23716 43120
rect 23204 42900 23256 42906
rect 23204 42842 23256 42848
rect 23020 42696 23072 42702
rect 23020 42638 23072 42644
rect 23768 42634 23796 43250
rect 23756 42628 23808 42634
rect 23756 42570 23808 42576
rect 22928 42560 22980 42566
rect 22928 42502 22980 42508
rect 22652 42356 22704 42362
rect 22652 42298 22704 42304
rect 23768 42226 23796 42570
rect 24044 42226 24072 43250
rect 23756 42220 23808 42226
rect 23756 42162 23808 42168
rect 24032 42220 24084 42226
rect 24032 42162 24084 42168
rect 24596 42158 24624 43318
rect 24584 42152 24636 42158
rect 24584 42094 24636 42100
rect 22008 42016 22060 42022
rect 22008 41958 22060 41964
rect 22744 42016 22796 42022
rect 22744 41958 22796 41964
rect 21192 41386 21312 41414
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 21284 7546 21312 41386
rect 22756 41274 22784 41958
rect 24780 41818 24808 43726
rect 25240 43314 25268 44338
rect 25228 43308 25280 43314
rect 25228 43250 25280 43256
rect 25240 42906 25268 43250
rect 25228 42900 25280 42906
rect 25228 42842 25280 42848
rect 25412 42696 25464 42702
rect 25412 42638 25464 42644
rect 25424 42294 25452 42638
rect 25412 42288 25464 42294
rect 25412 42230 25464 42236
rect 24768 41812 24820 41818
rect 24768 41754 24820 41760
rect 22744 41268 22796 41274
rect 22744 41210 22796 41216
rect 25976 41206 26004 44814
rect 26068 44402 26096 44950
rect 26252 44878 26280 45902
rect 26344 45354 26372 45902
rect 26436 45898 26464 46446
rect 26424 45892 26476 45898
rect 26476 45852 26556 45880
rect 26424 45834 26476 45840
rect 26424 45416 26476 45422
rect 26424 45358 26476 45364
rect 26332 45348 26384 45354
rect 26332 45290 26384 45296
rect 26240 44872 26292 44878
rect 26240 44814 26292 44820
rect 26344 44538 26372 45290
rect 26436 44878 26464 45358
rect 26424 44872 26476 44878
rect 26424 44814 26476 44820
rect 26332 44532 26384 44538
rect 26332 44474 26384 44480
rect 26056 44396 26108 44402
rect 26056 44338 26108 44344
rect 26068 43314 26096 44338
rect 26056 43308 26108 43314
rect 26056 43250 26108 43256
rect 26240 42900 26292 42906
rect 26240 42842 26292 42848
rect 26252 42362 26280 42842
rect 26240 42356 26292 42362
rect 26240 42298 26292 42304
rect 26252 41614 26280 42298
rect 26240 41608 26292 41614
rect 26240 41550 26292 41556
rect 26528 41274 26556 45852
rect 26620 45354 26648 49286
rect 26790 49200 26846 50000
rect 27158 49314 27214 50000
rect 26896 49286 27214 49314
rect 26804 46510 26832 49200
rect 26896 46986 26924 49286
rect 27158 49200 27214 49286
rect 27526 49200 27582 50000
rect 27894 49200 27950 50000
rect 28262 49200 28318 50000
rect 28630 49314 28686 50000
rect 28998 49314 29054 50000
rect 29366 49314 29422 50000
rect 28630 49286 28948 49314
rect 28630 49200 28686 49286
rect 26884 46980 26936 46986
rect 26884 46922 26936 46928
rect 27160 46980 27212 46986
rect 27160 46922 27212 46928
rect 27172 46646 27200 46922
rect 27160 46640 27212 46646
rect 27160 46582 27212 46588
rect 26976 46572 27028 46578
rect 26976 46514 27028 46520
rect 27068 46572 27120 46578
rect 27068 46514 27120 46520
rect 26792 46504 26844 46510
rect 26792 46446 26844 46452
rect 26988 45966 27016 46514
rect 27080 46170 27108 46514
rect 27068 46164 27120 46170
rect 27068 46106 27120 46112
rect 26976 45960 27028 45966
rect 26976 45902 27028 45908
rect 27540 45626 27568 49200
rect 27804 47116 27856 47122
rect 27804 47058 27856 47064
rect 27712 47048 27764 47054
rect 27712 46990 27764 46996
rect 27724 46170 27752 46990
rect 27816 46646 27844 47058
rect 27804 46640 27856 46646
rect 27804 46582 27856 46588
rect 27712 46164 27764 46170
rect 27712 46106 27764 46112
rect 27908 46034 27936 49200
rect 27896 46028 27948 46034
rect 27896 45970 27948 45976
rect 27620 45892 27672 45898
rect 27620 45834 27672 45840
rect 27528 45620 27580 45626
rect 27528 45562 27580 45568
rect 26608 45348 26660 45354
rect 26608 45290 26660 45296
rect 27252 45280 27304 45286
rect 27252 45222 27304 45228
rect 27160 44804 27212 44810
rect 27160 44746 27212 44752
rect 27172 43314 27200 44746
rect 27264 43926 27292 45222
rect 27632 44878 27660 45834
rect 27804 45824 27856 45830
rect 27804 45766 27856 45772
rect 27816 45286 27844 45766
rect 27988 45348 28040 45354
rect 27988 45290 28040 45296
rect 27804 45280 27856 45286
rect 27804 45222 27856 45228
rect 27620 44872 27672 44878
rect 27620 44814 27672 44820
rect 27632 44402 27660 44814
rect 27816 44538 27844 45222
rect 28000 44878 28028 45290
rect 27988 44872 28040 44878
rect 27988 44814 28040 44820
rect 27804 44532 27856 44538
rect 27804 44474 27856 44480
rect 27620 44396 27672 44402
rect 27620 44338 27672 44344
rect 27344 44328 27396 44334
rect 27344 44270 27396 44276
rect 27252 43920 27304 43926
rect 27252 43862 27304 43868
rect 27160 43308 27212 43314
rect 27160 43250 27212 43256
rect 27172 42634 27200 43250
rect 27264 43178 27292 43862
rect 27356 43790 27384 44270
rect 27816 43790 27844 44474
rect 28000 44470 28028 44814
rect 28172 44736 28224 44742
rect 28172 44678 28224 44684
rect 27988 44464 28040 44470
rect 27988 44406 28040 44412
rect 28184 44266 28212 44678
rect 28172 44260 28224 44266
rect 28172 44202 28224 44208
rect 28276 43994 28304 49200
rect 28920 47054 28948 49286
rect 28998 49286 29316 49314
rect 28998 49200 29054 49286
rect 28908 47048 28960 47054
rect 28908 46990 28960 46996
rect 29092 46572 29144 46578
rect 29092 46514 29144 46520
rect 28908 45960 28960 45966
rect 28908 45902 28960 45908
rect 28920 45490 28948 45902
rect 29000 45892 29052 45898
rect 29000 45834 29052 45840
rect 28908 45484 28960 45490
rect 28908 45426 28960 45432
rect 29012 45422 29040 45834
rect 28448 45416 28500 45422
rect 28448 45358 28500 45364
rect 29000 45416 29052 45422
rect 29000 45358 29052 45364
rect 28460 44402 28488 45358
rect 28448 44396 28500 44402
rect 28448 44338 28500 44344
rect 29012 44334 29040 45358
rect 29104 44470 29132 46514
rect 29288 45626 29316 49286
rect 29366 49286 29684 49314
rect 29366 49200 29422 49286
rect 29368 46912 29420 46918
rect 29368 46854 29420 46860
rect 29656 46866 29684 49286
rect 29734 49200 29790 50000
rect 30102 49200 30158 50000
rect 30470 49200 30526 50000
rect 30838 49314 30894 50000
rect 30576 49286 30894 49314
rect 29748 47002 29776 49200
rect 30012 47048 30064 47054
rect 29748 46974 29960 47002
rect 30012 46990 30064 46996
rect 29828 46912 29880 46918
rect 29656 46860 29828 46866
rect 29656 46854 29880 46860
rect 29380 46102 29408 46854
rect 29656 46838 29868 46854
rect 29644 46572 29696 46578
rect 29644 46514 29696 46520
rect 29656 46170 29684 46514
rect 29644 46164 29696 46170
rect 29644 46106 29696 46112
rect 29368 46096 29420 46102
rect 29368 46038 29420 46044
rect 29550 46064 29606 46073
rect 29380 45966 29408 46038
rect 29550 45999 29606 46008
rect 29368 45960 29420 45966
rect 29368 45902 29420 45908
rect 29276 45620 29328 45626
rect 29276 45562 29328 45568
rect 29564 45286 29592 45999
rect 29552 45280 29604 45286
rect 29552 45222 29604 45228
rect 29564 44878 29592 45222
rect 29656 44946 29684 46106
rect 29828 45960 29880 45966
rect 29828 45902 29880 45908
rect 29736 45416 29788 45422
rect 29736 45358 29788 45364
rect 29748 45014 29776 45358
rect 29736 45008 29788 45014
rect 29736 44950 29788 44956
rect 29644 44940 29696 44946
rect 29644 44882 29696 44888
rect 29552 44872 29604 44878
rect 29552 44814 29604 44820
rect 29092 44464 29144 44470
rect 29092 44406 29144 44412
rect 29748 44334 29776 44950
rect 29840 44402 29868 45902
rect 29932 45490 29960 46974
rect 30024 45490 30052 46990
rect 29920 45484 29972 45490
rect 29920 45426 29972 45432
rect 30012 45484 30064 45490
rect 30012 45426 30064 45432
rect 29828 44396 29880 44402
rect 29828 44338 29880 44344
rect 29000 44328 29052 44334
rect 29000 44270 29052 44276
rect 29736 44328 29788 44334
rect 29736 44270 29788 44276
rect 28264 43988 28316 43994
rect 28264 43930 28316 43936
rect 27344 43784 27396 43790
rect 27344 43726 27396 43732
rect 27620 43784 27672 43790
rect 27620 43726 27672 43732
rect 27804 43784 27856 43790
rect 27804 43726 27856 43732
rect 28080 43784 28132 43790
rect 28080 43726 28132 43732
rect 28172 43784 28224 43790
rect 28172 43726 28224 43732
rect 27632 43382 27660 43726
rect 27620 43376 27672 43382
rect 27620 43318 27672 43324
rect 27816 43314 27844 43726
rect 27988 43716 28040 43722
rect 27988 43658 28040 43664
rect 27804 43308 27856 43314
rect 27804 43250 27856 43256
rect 28000 43246 28028 43658
rect 27620 43240 27672 43246
rect 27620 43182 27672 43188
rect 27988 43240 28040 43246
rect 27988 43182 28040 43188
rect 27252 43172 27304 43178
rect 27252 43114 27304 43120
rect 27632 42702 27660 43182
rect 28000 42702 28028 43182
rect 28092 42770 28120 43726
rect 28184 43450 28212 43726
rect 28172 43444 28224 43450
rect 28172 43386 28224 43392
rect 28540 43308 28592 43314
rect 28540 43250 28592 43256
rect 28080 42764 28132 42770
rect 28080 42706 28132 42712
rect 27620 42696 27672 42702
rect 27620 42638 27672 42644
rect 27988 42696 28040 42702
rect 27988 42638 28040 42644
rect 28172 42696 28224 42702
rect 28172 42638 28224 42644
rect 27160 42628 27212 42634
rect 27160 42570 27212 42576
rect 26608 42016 26660 42022
rect 26608 41958 26660 41964
rect 26620 41614 26648 41958
rect 26608 41608 26660 41614
rect 26608 41550 26660 41556
rect 27632 41546 27660 42638
rect 28184 41818 28212 42638
rect 28172 41812 28224 41818
rect 28172 41754 28224 41760
rect 27620 41540 27672 41546
rect 27620 41482 27672 41488
rect 27344 41472 27396 41478
rect 27344 41414 27396 41420
rect 27356 41274 27384 41414
rect 28552 41274 28580 43250
rect 29748 43246 29776 44270
rect 30024 43314 30052 45426
rect 30116 43994 30144 49200
rect 30288 47116 30340 47122
rect 30288 47058 30340 47064
rect 30300 45966 30328 47058
rect 30380 46980 30432 46986
rect 30380 46922 30432 46928
rect 30392 46714 30420 46922
rect 30484 46889 30512 49200
rect 30470 46880 30526 46889
rect 30470 46815 30526 46824
rect 30380 46708 30432 46714
rect 30380 46650 30432 46656
rect 30472 46572 30524 46578
rect 30472 46514 30524 46520
rect 30288 45960 30340 45966
rect 30288 45902 30340 45908
rect 30196 45892 30248 45898
rect 30196 45834 30248 45840
rect 30104 43988 30156 43994
rect 30104 43930 30156 43936
rect 30012 43308 30064 43314
rect 30012 43250 30064 43256
rect 29736 43240 29788 43246
rect 29736 43182 29788 43188
rect 29644 42832 29696 42838
rect 29644 42774 29696 42780
rect 29460 42628 29512 42634
rect 29460 42570 29512 42576
rect 29472 42226 29500 42570
rect 29460 42220 29512 42226
rect 29460 42162 29512 42168
rect 26240 41268 26292 41274
rect 26240 41210 26292 41216
rect 26516 41268 26568 41274
rect 26516 41210 26568 41216
rect 27344 41268 27396 41274
rect 27344 41210 27396 41216
rect 28540 41268 28592 41274
rect 28540 41210 28592 41216
rect 25964 41200 26016 41206
rect 25964 41142 26016 41148
rect 26252 41138 26280 41210
rect 26240 41132 26292 41138
rect 26240 41074 26292 41080
rect 29656 40934 29684 42774
rect 29748 42770 29776 43182
rect 30024 42838 30052 43250
rect 30012 42832 30064 42838
rect 30012 42774 30064 42780
rect 29736 42764 29788 42770
rect 29736 42706 29788 42712
rect 30208 42634 30236 45834
rect 30300 44946 30328 45902
rect 30380 45348 30432 45354
rect 30380 45290 30432 45296
rect 30288 44940 30340 44946
rect 30288 44882 30340 44888
rect 30392 43382 30420 45290
rect 30380 43376 30432 43382
rect 30380 43318 30432 43324
rect 30392 42702 30420 43318
rect 30380 42696 30432 42702
rect 30380 42638 30432 42644
rect 30196 42628 30248 42634
rect 30196 42570 30248 42576
rect 30208 41206 30236 42570
rect 30484 41546 30512 46514
rect 30576 43926 30604 49286
rect 30838 49200 30894 49286
rect 31206 49314 31262 50000
rect 31206 49286 31524 49314
rect 31206 49200 31262 49286
rect 31208 47116 31260 47122
rect 31208 47058 31260 47064
rect 30840 47048 30892 47054
rect 30892 47008 30972 47036
rect 30840 46990 30892 46996
rect 30944 46510 30972 47008
rect 31220 46968 31248 47058
rect 31300 47048 31352 47054
rect 31300 46990 31352 46996
rect 31128 46940 31248 46968
rect 31128 46510 31156 46940
rect 31312 46578 31340 46990
rect 31300 46572 31352 46578
rect 31300 46514 31352 46520
rect 30932 46504 30984 46510
rect 30932 46446 30984 46452
rect 31116 46504 31168 46510
rect 31116 46446 31168 46452
rect 30944 46102 30972 46446
rect 30932 46096 30984 46102
rect 30932 46038 30984 46044
rect 31024 45484 31076 45490
rect 31024 45426 31076 45432
rect 30564 43920 30616 43926
rect 30564 43862 30616 43868
rect 30576 43314 30604 43862
rect 30564 43308 30616 43314
rect 30564 43250 30616 43256
rect 30576 42362 30604 43250
rect 30656 42560 30708 42566
rect 30656 42502 30708 42508
rect 30668 42362 30696 42502
rect 31036 42362 31064 45426
rect 31128 43994 31156 46446
rect 31312 46170 31340 46514
rect 31300 46164 31352 46170
rect 31300 46106 31352 46112
rect 31496 45830 31524 49286
rect 31574 49200 31630 50000
rect 31942 49314 31998 50000
rect 31942 49286 32260 49314
rect 31942 49200 31998 49286
rect 31588 46646 31616 49200
rect 32036 46980 32088 46986
rect 32036 46922 32088 46928
rect 31576 46640 31628 46646
rect 31576 46582 31628 46588
rect 32048 45966 32076 46922
rect 32036 45960 32088 45966
rect 32036 45902 32088 45908
rect 31944 45892 31996 45898
rect 31944 45834 31996 45840
rect 31484 45824 31536 45830
rect 31484 45766 31536 45772
rect 31956 44878 31984 45834
rect 31944 44872 31996 44878
rect 31944 44814 31996 44820
rect 32036 44872 32088 44878
rect 32036 44814 32088 44820
rect 31956 44402 31984 44814
rect 31944 44396 31996 44402
rect 31944 44338 31996 44344
rect 31852 44328 31904 44334
rect 31588 44266 31800 44282
rect 31852 44270 31904 44276
rect 31576 44260 31800 44266
rect 31628 44254 31800 44260
rect 31576 44202 31628 44208
rect 31772 43994 31800 44254
rect 31116 43988 31168 43994
rect 31116 43930 31168 43936
rect 31760 43988 31812 43994
rect 31760 43930 31812 43936
rect 31864 43790 31892 44270
rect 32048 44198 32076 44814
rect 32036 44192 32088 44198
rect 32036 44134 32088 44140
rect 31852 43784 31904 43790
rect 31852 43726 31904 43732
rect 31300 43172 31352 43178
rect 31300 43114 31352 43120
rect 30564 42356 30616 42362
rect 30564 42298 30616 42304
rect 30656 42356 30708 42362
rect 30656 42298 30708 42304
rect 31024 42356 31076 42362
rect 31024 42298 31076 42304
rect 30668 42226 30696 42298
rect 30656 42220 30708 42226
rect 30656 42162 30708 42168
rect 31312 41818 31340 43114
rect 32232 42226 32260 49286
rect 32310 49200 32366 50000
rect 32678 49200 32734 50000
rect 33046 49200 33102 50000
rect 33414 49314 33470 50000
rect 33782 49314 33838 50000
rect 34150 49314 34206 50000
rect 34518 49314 34574 50000
rect 34886 49314 34942 50000
rect 35254 49314 35310 50000
rect 33414 49286 33732 49314
rect 33414 49200 33470 49286
rect 32324 46442 32352 49200
rect 32692 46714 32720 49200
rect 32680 46708 32732 46714
rect 32680 46650 32732 46656
rect 32312 46436 32364 46442
rect 32312 46378 32364 46384
rect 33060 46374 33088 49200
rect 33704 47410 33732 49286
rect 33782 49286 34100 49314
rect 33782 49200 33838 49286
rect 34072 47546 34100 49286
rect 34150 49286 34468 49314
rect 34150 49200 34206 49286
rect 34072 47518 34376 47546
rect 33704 47382 34284 47410
rect 33876 47184 33928 47190
rect 33876 47126 33928 47132
rect 33692 47048 33744 47054
rect 33692 46990 33744 46996
rect 33140 46980 33192 46986
rect 33140 46922 33192 46928
rect 33152 46578 33180 46922
rect 33598 46744 33654 46753
rect 33598 46679 33654 46688
rect 33612 46646 33640 46679
rect 33508 46640 33560 46646
rect 33508 46582 33560 46588
rect 33600 46640 33652 46646
rect 33600 46582 33652 46588
rect 33140 46572 33192 46578
rect 33140 46514 33192 46520
rect 33232 46572 33284 46578
rect 33232 46514 33284 46520
rect 33048 46368 33100 46374
rect 33048 46310 33100 46316
rect 33152 46034 33180 46514
rect 33244 46170 33272 46514
rect 33232 46164 33284 46170
rect 33232 46106 33284 46112
rect 33520 46034 33548 46582
rect 33140 46028 33192 46034
rect 33140 45970 33192 45976
rect 33508 46028 33560 46034
rect 33508 45970 33560 45976
rect 33704 45966 33732 46990
rect 33888 45966 33916 47126
rect 34152 46708 34204 46714
rect 34152 46650 34204 46656
rect 33416 45960 33468 45966
rect 33416 45902 33468 45908
rect 33692 45960 33744 45966
rect 33692 45902 33744 45908
rect 33876 45960 33928 45966
rect 33928 45920 34008 45948
rect 33876 45902 33928 45908
rect 33428 45490 33456 45902
rect 33048 45484 33100 45490
rect 33048 45426 33100 45432
rect 33416 45484 33468 45490
rect 33416 45426 33468 45432
rect 32312 44872 32364 44878
rect 32312 44814 32364 44820
rect 32324 43994 32352 44814
rect 33060 44146 33088 45426
rect 33416 44940 33468 44946
rect 33416 44882 33468 44888
rect 33140 44804 33192 44810
rect 33140 44746 33192 44752
rect 33152 44334 33180 44746
rect 33428 44470 33456 44882
rect 33980 44878 34008 45920
rect 34060 45892 34112 45898
rect 34060 45834 34112 45840
rect 34072 45422 34100 45834
rect 34060 45416 34112 45422
rect 34060 45358 34112 45364
rect 34072 44946 34100 45358
rect 34164 45082 34192 46650
rect 34152 45076 34204 45082
rect 34152 45018 34204 45024
rect 34060 44940 34112 44946
rect 34060 44882 34112 44888
rect 33968 44872 34020 44878
rect 33968 44814 34020 44820
rect 33416 44464 33468 44470
rect 33416 44406 33468 44412
rect 33140 44328 33192 44334
rect 33140 44270 33192 44276
rect 33060 44118 33180 44146
rect 32312 43988 32364 43994
rect 32312 43930 32364 43936
rect 32772 43784 32824 43790
rect 32772 43726 32824 43732
rect 32784 43382 32812 43726
rect 32772 43376 32824 43382
rect 32772 43318 32824 43324
rect 33152 42770 33180 44118
rect 33140 42764 33192 42770
rect 33140 42706 33192 42712
rect 32404 42696 32456 42702
rect 32404 42638 32456 42644
rect 32220 42220 32272 42226
rect 32220 42162 32272 42168
rect 31300 41812 31352 41818
rect 31300 41754 31352 41760
rect 30472 41540 30524 41546
rect 30472 41482 30524 41488
rect 30840 41540 30892 41546
rect 30840 41482 30892 41488
rect 30196 41200 30248 41206
rect 30196 41142 30248 41148
rect 29644 40928 29696 40934
rect 29644 40870 29696 40876
rect 29656 40730 29684 40870
rect 29644 40724 29696 40730
rect 29644 40666 29696 40672
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 24032 7880 24084 7886
rect 24032 7822 24084 7828
rect 24952 7880 25004 7886
rect 24952 7822 25004 7828
rect 26056 7880 26108 7886
rect 26056 7822 26108 7828
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 21284 6798 21312 7482
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 22112 6662 22140 7346
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 22284 6656 22336 6662
rect 22284 6598 22336 6604
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 18236 5160 18288 5166
rect 18236 5102 18288 5108
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 18248 4826 18276 5102
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 19352 4622 19380 6598
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 20548 5914 20576 6326
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20916 5710 20944 6598
rect 21088 6248 21140 6254
rect 21088 6190 21140 6196
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20904 5704 20956 5710
rect 20904 5646 20956 5652
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 20088 5302 20116 5510
rect 20076 5296 20128 5302
rect 20076 5238 20128 5244
rect 20364 4622 20392 5646
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 4172 2938 4200 3470
rect 4080 2910 4200 2938
rect 4896 2916 4948 2922
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2608 800 2636 2382
rect 3160 800 3188 2790
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 3528 800 3556 2450
rect 3896 800 3924 2790
rect 4080 2564 4108 2910
rect 4896 2858 4948 2864
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4080 2536 4292 2564
rect 4264 800 4292 2536
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4632 800 4660 2382
rect 4908 800 4936 2858
rect 5184 800 5212 3470
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5460 800 5488 2926
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5736 800 5764 2382
rect 6012 800 6040 3470
rect 6276 2916 6328 2922
rect 6276 2858 6328 2864
rect 6288 800 6316 2858
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6564 800 6592 2790
rect 6840 800 6868 3470
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7116 800 7144 2518
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 7392 800 7420 2314
rect 7668 800 7696 3470
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7944 800 7972 2926
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8220 800 8248 2450
rect 8496 800 8524 3470
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8772 800 8800 2858
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 9048 800 9076 2790
rect 9324 800 9352 3470
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9588 2576 9640 2582
rect 9588 2518 9640 2524
rect 9600 800 9628 2518
rect 9876 800 9904 2926
rect 10152 800 10180 3470
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 10416 2508 10468 2514
rect 10416 2450 10468 2456
rect 10428 800 10456 2450
rect 10704 800 10732 2790
rect 10980 800 11008 3470
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11256 800 11284 2858
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 11532 800 11560 2518
rect 11808 800 11836 3470
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12084 800 12112 2790
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12268 800 12296 2382
rect 12544 800 12572 3470
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 12820 800 12848 2450
rect 13096 800 13124 3470
rect 13360 2916 13412 2922
rect 13360 2858 13412 2864
rect 13372 800 13400 2858
rect 13648 800 13676 3470
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13924 800 13952 2790
rect 14188 2576 14240 2582
rect 14188 2518 14240 2524
rect 14200 800 14228 2518
rect 14476 800 14504 2858
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 14752 800 14780 2450
rect 15028 800 15056 3470
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 15304 800 15332 2926
rect 15844 2848 15896 2854
rect 15844 2790 15896 2796
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15580 800 15608 2382
rect 15856 800 15884 2790
rect 16132 800 16160 3878
rect 16856 3664 16908 3670
rect 16856 3606 16908 3612
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16408 800 16436 3470
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 16684 800 16712 2450
rect 16868 1850 16896 3606
rect 16868 1822 16988 1850
rect 16960 800 16988 1822
rect 17236 800 17264 3878
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17512 800 17540 2926
rect 17788 800 17816 3538
rect 18052 2916 18104 2922
rect 18052 2858 18104 2864
rect 18064 800 18092 2858
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 18340 800 18368 2314
rect 18616 800 18644 3946
rect 19352 3670 19380 4558
rect 20364 4486 20392 4558
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 20364 4146 20392 4422
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19156 3664 19208 3670
rect 19156 3606 19208 3612
rect 19340 3664 19392 3670
rect 19340 3606 19392 3612
rect 18880 3460 18932 3466
rect 18880 3402 18932 3408
rect 18892 3058 18920 3402
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 18892 800 18920 2450
rect 19168 800 19196 3606
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19352 2650 19380 2926
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19444 800 19472 3878
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 1442 20024 2790
rect 19720 1414 20024 1442
rect 19720 800 19748 1414
rect 20088 1306 20116 3674
rect 20168 3460 20220 3466
rect 20168 3402 20220 3408
rect 20180 3194 20208 3402
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 20364 3058 20392 4082
rect 20536 3120 20588 3126
rect 20536 3062 20588 3068
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 20260 2576 20312 2582
rect 20260 2518 20312 2524
rect 19996 1278 20116 1306
rect 19996 800 20024 1278
rect 20272 800 20300 2518
rect 20364 2378 20392 2994
rect 20352 2372 20404 2378
rect 20352 2314 20404 2320
rect 20548 800 20576 3062
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 20824 800 20852 2382
rect 21100 800 21128 6190
rect 21560 5710 21588 6598
rect 22296 5778 22324 6598
rect 22480 6254 22508 7142
rect 23032 6866 23060 7822
rect 23112 7200 23164 7206
rect 23112 7142 23164 7148
rect 23020 6860 23072 6866
rect 23020 6802 23072 6808
rect 23124 6730 23152 7142
rect 23848 6860 23900 6866
rect 23848 6802 23900 6808
rect 23112 6724 23164 6730
rect 23112 6666 23164 6672
rect 23388 6724 23440 6730
rect 23388 6666 23440 6672
rect 22560 6384 22612 6390
rect 22560 6326 22612 6332
rect 22468 6248 22520 6254
rect 22468 6190 22520 6196
rect 22572 5914 22600 6326
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 23400 5710 23428 6666
rect 23572 6248 23624 6254
rect 23572 6190 23624 6196
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 22836 5704 22888 5710
rect 22836 5646 22888 5652
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 21180 5024 21232 5030
rect 21180 4966 21232 4972
rect 21192 4690 21220 4966
rect 21180 4684 21232 4690
rect 21180 4626 21232 4632
rect 21456 4140 21508 4146
rect 21456 4082 21508 4088
rect 21272 3936 21324 3942
rect 21468 3924 21496 4082
rect 21324 3896 21496 3924
rect 21272 3878 21324 3884
rect 21560 3534 21588 5646
rect 22652 5636 22704 5642
rect 22652 5578 22704 5584
rect 22664 5302 22692 5578
rect 22652 5296 22704 5302
rect 22652 5238 22704 5244
rect 21640 5160 21692 5166
rect 21640 5102 21692 5108
rect 22560 5160 22612 5166
rect 22560 5102 22612 5108
rect 21548 3528 21600 3534
rect 21548 3470 21600 3476
rect 21364 3460 21416 3466
rect 21364 3402 21416 3408
rect 21376 800 21404 3402
rect 21560 3058 21588 3470
rect 21548 3052 21600 3058
rect 21548 2994 21600 3000
rect 21652 800 21680 5102
rect 22572 4826 22600 5102
rect 22560 4820 22612 4826
rect 22560 4762 22612 4768
rect 21824 4684 21876 4690
rect 21824 4626 21876 4632
rect 21836 2258 21864 4626
rect 22848 4622 22876 5646
rect 23204 5160 23256 5166
rect 23204 5102 23256 5108
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 22848 4282 22876 4558
rect 22836 4276 22888 4282
rect 22836 4218 22888 4224
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 22204 2650 22232 3062
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 21836 2230 21956 2258
rect 21928 800 21956 2230
rect 22296 2122 22324 4014
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22468 2984 22520 2990
rect 22468 2926 22520 2932
rect 22204 2094 22324 2122
rect 22204 800 22232 2094
rect 22480 800 22508 2926
rect 22756 800 22784 3538
rect 22836 2848 22888 2854
rect 22836 2790 22888 2796
rect 22848 2378 22876 2790
rect 23020 2508 23072 2514
rect 23020 2450 23072 2456
rect 22836 2372 22888 2378
rect 22836 2314 22888 2320
rect 23032 800 23060 2450
rect 23216 2258 23244 5102
rect 23480 4548 23532 4554
rect 23480 4490 23532 4496
rect 23492 4214 23520 4490
rect 23480 4208 23532 4214
rect 23480 4150 23532 4156
rect 23216 2230 23336 2258
rect 23308 800 23336 2230
rect 23584 800 23612 6190
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23768 3126 23796 3878
rect 23756 3120 23808 3126
rect 23756 3062 23808 3068
rect 23860 800 23888 6802
rect 24044 6390 24072 7822
rect 24964 7478 24992 7822
rect 25412 7744 25464 7750
rect 25412 7686 25464 7692
rect 24860 7472 24912 7478
rect 24860 7414 24912 7420
rect 24952 7472 25004 7478
rect 24952 7414 25004 7420
rect 24872 7002 24900 7414
rect 25228 7336 25280 7342
rect 25228 7278 25280 7284
rect 24860 6996 24912 7002
rect 24860 6938 24912 6944
rect 24032 6384 24084 6390
rect 24032 6326 24084 6332
rect 24124 6384 24176 6390
rect 24124 6326 24176 6332
rect 24136 5914 24164 6326
rect 24952 6248 25004 6254
rect 24952 6190 25004 6196
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 24308 5636 24360 5642
rect 24308 5578 24360 5584
rect 24320 5302 24348 5578
rect 24308 5296 24360 5302
rect 24308 5238 24360 5244
rect 24860 5160 24912 5166
rect 24860 5102 24912 5108
rect 24124 4072 24176 4078
rect 24124 4014 24176 4020
rect 24136 800 24164 4014
rect 24400 2984 24452 2990
rect 24400 2926 24452 2932
rect 24584 2984 24636 2990
rect 24584 2926 24636 2932
rect 24412 800 24440 2926
rect 24596 2310 24624 2926
rect 24872 2802 24900 5102
rect 24688 2774 24900 2802
rect 24584 2304 24636 2310
rect 24584 2246 24636 2252
rect 24688 800 24716 2774
rect 24964 800 24992 6190
rect 25044 4548 25096 4554
rect 25044 4490 25096 4496
rect 25056 2378 25084 4490
rect 25044 2372 25096 2378
rect 25044 2314 25096 2320
rect 25240 800 25268 7278
rect 25424 6798 25452 7686
rect 25688 7472 25740 7478
rect 25688 7414 25740 7420
rect 25700 7002 25728 7414
rect 26068 7342 26096 7822
rect 26148 7812 26200 7818
rect 26148 7754 26200 7760
rect 26056 7336 26108 7342
rect 26056 7278 26108 7284
rect 25688 6996 25740 7002
rect 25688 6938 25740 6944
rect 25412 6792 25464 6798
rect 25412 6734 25464 6740
rect 25424 5710 25452 6734
rect 26160 6662 26188 7754
rect 26608 7336 26660 7342
rect 26608 7278 26660 7284
rect 26240 7200 26292 7206
rect 26240 7142 26292 7148
rect 26148 6656 26200 6662
rect 26148 6598 26200 6604
rect 25688 6384 25740 6390
rect 25688 6326 25740 6332
rect 25700 5914 25728 6326
rect 25688 5908 25740 5914
rect 25688 5850 25740 5856
rect 26160 5778 26188 6598
rect 26252 6254 26280 7142
rect 26516 6316 26568 6322
rect 26516 6258 26568 6264
rect 26240 6248 26292 6254
rect 26240 6190 26292 6196
rect 26332 6180 26384 6186
rect 26332 6122 26384 6128
rect 26148 5772 26200 5778
rect 26148 5714 26200 5720
rect 25412 5704 25464 5710
rect 25412 5646 25464 5652
rect 25424 5250 25452 5646
rect 25424 5222 25544 5250
rect 25516 4690 25544 5222
rect 25504 4684 25556 4690
rect 25504 4626 25556 4632
rect 25964 4684 26016 4690
rect 25964 4626 26016 4632
rect 25412 4548 25464 4554
rect 25412 4490 25464 4496
rect 25424 4282 25452 4490
rect 25412 4276 25464 4282
rect 25412 4218 25464 4224
rect 25516 4146 25544 4626
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 25516 3534 25544 4082
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 25412 3392 25464 3398
rect 25412 3334 25464 3340
rect 25424 3126 25452 3334
rect 25412 3120 25464 3126
rect 25412 3062 25464 3068
rect 25780 2984 25832 2990
rect 25780 2926 25832 2932
rect 25504 2508 25556 2514
rect 25504 2450 25556 2456
rect 25516 800 25544 2450
rect 25792 800 25820 2926
rect 25976 2394 26004 4626
rect 25976 2366 26096 2394
rect 26068 800 26096 2366
rect 26344 800 26372 6122
rect 26528 5914 26556 6258
rect 26516 5908 26568 5914
rect 26516 5850 26568 5856
rect 26528 5234 26556 5850
rect 26516 5228 26568 5234
rect 26516 5170 26568 5176
rect 26424 4480 26476 4486
rect 26424 4422 26476 4428
rect 26436 2650 26464 4422
rect 26528 4146 26556 5170
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 26528 3534 26556 4082
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26424 2644 26476 2650
rect 26424 2586 26476 2592
rect 26620 800 26648 7278
rect 27712 7200 27764 7206
rect 27712 7142 27764 7148
rect 27724 6866 27752 7142
rect 27712 6860 27764 6866
rect 27712 6802 27764 6808
rect 27988 6860 28040 6866
rect 27988 6802 28040 6808
rect 27804 6724 27856 6730
rect 27804 6666 27856 6672
rect 27816 6458 27844 6666
rect 27804 6452 27856 6458
rect 27804 6394 27856 6400
rect 27712 5772 27764 5778
rect 27712 5714 27764 5720
rect 27252 5160 27304 5166
rect 27252 5102 27304 5108
rect 27620 5160 27672 5166
rect 27620 5102 27672 5108
rect 27264 4826 27292 5102
rect 27252 4820 27304 4826
rect 27252 4762 27304 4768
rect 26884 4072 26936 4078
rect 26884 4014 26936 4020
rect 26896 800 26924 4014
rect 27160 2984 27212 2990
rect 27160 2926 27212 2932
rect 27172 800 27200 2926
rect 27632 2802 27660 5102
rect 27448 2774 27660 2802
rect 27448 800 27476 2774
rect 27724 800 27752 5714
rect 28000 800 28028 6802
rect 29000 6656 29052 6662
rect 29000 6598 29052 6604
rect 28172 6112 28224 6118
rect 28172 6054 28224 6060
rect 28184 5642 28212 6054
rect 29012 5710 29040 6598
rect 29736 6112 29788 6118
rect 29736 6054 29788 6060
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 28172 5636 28224 5642
rect 28172 5578 28224 5584
rect 28264 5636 28316 5642
rect 28264 5578 28316 5584
rect 28276 4826 28304 5578
rect 28816 5160 28868 5166
rect 28816 5102 28868 5108
rect 28264 4820 28316 4826
rect 28264 4762 28316 4768
rect 28724 3936 28776 3942
rect 28724 3878 28776 3884
rect 28540 3596 28592 3602
rect 28540 3538 28592 3544
rect 28080 3392 28132 3398
rect 28080 3334 28132 3340
rect 28092 3126 28120 3334
rect 28080 3120 28132 3126
rect 28080 3062 28132 3068
rect 28264 2508 28316 2514
rect 28264 2450 28316 2456
rect 28276 800 28304 2450
rect 28552 800 28580 3538
rect 28736 3466 28764 3878
rect 28724 3460 28776 3466
rect 28724 3402 28776 3408
rect 28828 800 28856 5102
rect 29012 4842 29040 5646
rect 29644 5636 29696 5642
rect 29644 5578 29696 5584
rect 29656 5302 29684 5578
rect 29748 5302 29776 6054
rect 29644 5296 29696 5302
rect 29644 5238 29696 5244
rect 29736 5296 29788 5302
rect 29736 5238 29788 5244
rect 29012 4814 29224 4842
rect 29000 4684 29052 4690
rect 29052 4644 29132 4672
rect 29000 4626 29052 4632
rect 29104 800 29132 4644
rect 29196 4570 29224 4814
rect 29276 4616 29328 4622
rect 29196 4564 29276 4570
rect 29196 4558 29328 4564
rect 30104 4616 30156 4622
rect 30104 4558 30156 4564
rect 29196 4542 29316 4558
rect 29196 4146 29224 4542
rect 29184 4140 29236 4146
rect 29184 4082 29236 4088
rect 29736 3528 29788 3534
rect 29736 3470 29788 3476
rect 29920 3528 29972 3534
rect 29920 3470 29972 3476
rect 29644 3460 29696 3466
rect 29644 3402 29696 3408
rect 29184 2984 29236 2990
rect 29184 2926 29236 2932
rect 29368 2984 29420 2990
rect 29368 2926 29420 2932
rect 29196 2650 29224 2926
rect 29184 2644 29236 2650
rect 29184 2586 29236 2592
rect 29380 800 29408 2926
rect 29656 800 29684 3402
rect 29748 2514 29776 3470
rect 29736 2508 29788 2514
rect 29736 2450 29788 2456
rect 29932 800 29960 3470
rect 30116 3058 30144 4558
rect 30196 3936 30248 3942
rect 30196 3878 30248 3884
rect 30208 3602 30236 3878
rect 30196 3596 30248 3602
rect 30196 3538 30248 3544
rect 30472 3528 30524 3534
rect 30472 3470 30524 3476
rect 30104 3052 30156 3058
rect 30104 2994 30156 3000
rect 30116 2446 30144 2994
rect 30196 2848 30248 2854
rect 30196 2790 30248 2796
rect 30104 2440 30156 2446
rect 30104 2382 30156 2388
rect 30208 800 30236 2790
rect 30484 800 30512 3470
rect 30852 3466 30880 41482
rect 32416 41274 32444 42638
rect 33152 41750 33180 42706
rect 33428 42702 33456 44406
rect 33692 44328 33744 44334
rect 33692 44270 33744 44276
rect 33704 43858 33732 44270
rect 33692 43852 33744 43858
rect 33692 43794 33744 43800
rect 33784 43784 33836 43790
rect 33784 43726 33836 43732
rect 33796 43178 33824 43726
rect 33784 43172 33836 43178
rect 33784 43114 33836 43120
rect 33796 42770 33824 43114
rect 33784 42764 33836 42770
rect 33784 42706 33836 42712
rect 33416 42696 33468 42702
rect 33416 42638 33468 42644
rect 33980 42362 34008 44814
rect 34152 44192 34204 44198
rect 34152 44134 34204 44140
rect 34164 43790 34192 44134
rect 34152 43784 34204 43790
rect 34152 43726 34204 43732
rect 34164 43382 34192 43726
rect 34152 43376 34204 43382
rect 34152 43318 34204 43324
rect 34256 43314 34284 47382
rect 34348 46481 34376 47518
rect 34440 47138 34468 49286
rect 34518 49286 34744 49314
rect 34518 49200 34574 49286
rect 34440 47110 34560 47138
rect 34428 46980 34480 46986
rect 34428 46922 34480 46928
rect 34440 46578 34468 46922
rect 34428 46572 34480 46578
rect 34428 46514 34480 46520
rect 34334 46472 34390 46481
rect 34532 46458 34560 47110
rect 34612 46572 34664 46578
rect 34612 46514 34664 46520
rect 34334 46407 34390 46416
rect 34440 46430 34560 46458
rect 34336 46164 34388 46170
rect 34336 46106 34388 46112
rect 34348 44402 34376 46106
rect 34440 45898 34468 46430
rect 34428 45892 34480 45898
rect 34428 45834 34480 45840
rect 34624 44742 34652 46514
rect 34612 44736 34664 44742
rect 34612 44678 34664 44684
rect 34428 44464 34480 44470
rect 34428 44406 34480 44412
rect 34336 44396 34388 44402
rect 34336 44338 34388 44344
rect 34348 43738 34376 44338
rect 34440 44198 34468 44406
rect 34612 44396 34664 44402
rect 34612 44338 34664 44344
rect 34428 44192 34480 44198
rect 34428 44134 34480 44140
rect 34520 43784 34572 43790
rect 34348 43722 34468 43738
rect 34520 43726 34572 43732
rect 34348 43716 34480 43722
rect 34348 43710 34428 43716
rect 34244 43308 34296 43314
rect 34244 43250 34296 43256
rect 34348 42702 34376 43710
rect 34428 43658 34480 43664
rect 34532 43246 34560 43726
rect 34624 43654 34652 44338
rect 34612 43648 34664 43654
rect 34612 43590 34664 43596
rect 34520 43240 34572 43246
rect 34520 43182 34572 43188
rect 34624 43110 34652 43590
rect 34612 43104 34664 43110
rect 34612 43046 34664 43052
rect 34624 42770 34652 43046
rect 34716 42770 34744 49286
rect 34886 49286 35204 49314
rect 34886 49200 34942 49286
rect 35176 47546 35204 49286
rect 35254 49286 35572 49314
rect 35254 49200 35310 49286
rect 35176 47518 35480 47546
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 35348 46572 35400 46578
rect 35348 46514 35400 46520
rect 34796 46504 34848 46510
rect 34796 46446 34848 46452
rect 34808 45558 34836 46446
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34796 45552 34848 45558
rect 34796 45494 34848 45500
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 35360 45014 35388 46514
rect 34980 45008 35032 45014
rect 34980 44950 35032 44956
rect 35348 45008 35400 45014
rect 35348 44950 35400 44956
rect 34992 44470 35020 44950
rect 34980 44464 35032 44470
rect 34980 44406 35032 44412
rect 34796 44328 34848 44334
rect 34796 44270 34848 44276
rect 34808 43790 34836 44270
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34796 43784 34848 43790
rect 34796 43726 34848 43732
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 35452 42770 35480 47518
rect 35544 47054 35572 49286
rect 35622 49200 35678 50000
rect 35990 49200 36046 50000
rect 36358 49200 36414 50000
rect 36726 49200 36782 50000
rect 37094 49314 37150 50000
rect 37462 49314 37518 50000
rect 37094 49286 37228 49314
rect 37094 49200 37150 49286
rect 35532 47048 35584 47054
rect 35532 46990 35584 46996
rect 35544 46918 35572 46990
rect 35532 46912 35584 46918
rect 35532 46854 35584 46860
rect 35530 46608 35586 46617
rect 35530 46543 35532 46552
rect 35584 46543 35586 46552
rect 35532 46514 35584 46520
rect 35636 46374 35664 49200
rect 36004 46918 36032 49200
rect 36372 47190 36400 49200
rect 36360 47184 36412 47190
rect 36360 47126 36412 47132
rect 36360 47048 36412 47054
rect 36360 46990 36412 46996
rect 35716 46912 35768 46918
rect 35716 46854 35768 46860
rect 35992 46912 36044 46918
rect 36372 46889 36400 46990
rect 36636 46980 36688 46986
rect 36636 46922 36688 46928
rect 35992 46854 36044 46860
rect 36358 46880 36414 46889
rect 35624 46368 35676 46374
rect 35624 46310 35676 46316
rect 35728 46170 35756 46854
rect 36358 46815 36414 46824
rect 36648 46730 36676 46922
rect 36740 46889 36768 49200
rect 36820 47184 36872 47190
rect 36820 47126 36872 47132
rect 36726 46880 36782 46889
rect 36726 46815 36782 46824
rect 36648 46702 36768 46730
rect 36360 46504 36412 46510
rect 36360 46446 36412 46452
rect 36636 46504 36688 46510
rect 36636 46446 36688 46452
rect 36268 46436 36320 46442
rect 36268 46378 36320 46384
rect 35716 46164 35768 46170
rect 35716 46106 35768 46112
rect 36280 45626 36308 46378
rect 36372 46170 36400 46446
rect 36360 46164 36412 46170
rect 36360 46106 36412 46112
rect 36268 45620 36320 45626
rect 36268 45562 36320 45568
rect 36648 45558 36676 46446
rect 35624 45552 35676 45558
rect 35624 45494 35676 45500
rect 36636 45552 36688 45558
rect 36636 45494 36688 45500
rect 35532 45416 35584 45422
rect 35532 45358 35584 45364
rect 35544 44878 35572 45358
rect 35532 44872 35584 44878
rect 35532 44814 35584 44820
rect 35544 43722 35572 44814
rect 35636 44402 35664 45494
rect 36740 45490 36768 46702
rect 36832 46646 36860 47126
rect 37096 46912 37148 46918
rect 37096 46854 37148 46860
rect 36820 46640 36872 46646
rect 36820 46582 36872 46588
rect 36912 46504 36964 46510
rect 36912 46446 36964 46452
rect 36924 45966 36952 46446
rect 36912 45960 36964 45966
rect 36912 45902 36964 45908
rect 37108 45665 37136 46854
rect 37200 46753 37228 49286
rect 37292 49286 37518 49314
rect 37186 46744 37242 46753
rect 37186 46679 37242 46688
rect 37292 45778 37320 49286
rect 37462 49200 37518 49286
rect 37830 49200 37886 50000
rect 38198 49200 38254 50000
rect 38566 49200 38622 50000
rect 38934 49200 38990 50000
rect 39302 49200 39358 50000
rect 39670 49314 39726 50000
rect 39408 49286 39726 49314
rect 37648 47116 37700 47122
rect 37648 47058 37700 47064
rect 37464 47048 37516 47054
rect 37464 46990 37516 46996
rect 37476 46714 37504 46990
rect 37464 46708 37516 46714
rect 37464 46650 37516 46656
rect 37372 46436 37424 46442
rect 37372 46378 37424 46384
rect 37200 45750 37320 45778
rect 37094 45656 37150 45665
rect 37094 45591 37150 45600
rect 36728 45484 36780 45490
rect 36728 45426 36780 45432
rect 35716 45416 35768 45422
rect 35716 45358 35768 45364
rect 36268 45416 36320 45422
rect 36268 45358 36320 45364
rect 35728 44878 35756 45358
rect 36280 44946 36308 45358
rect 36268 44940 36320 44946
rect 36320 44900 36400 44928
rect 36268 44882 36320 44888
rect 35716 44872 35768 44878
rect 35716 44814 35768 44820
rect 35624 44396 35676 44402
rect 35624 44338 35676 44344
rect 35728 44334 35756 44814
rect 36176 44736 36228 44742
rect 36176 44678 36228 44684
rect 36188 44402 36216 44678
rect 36176 44396 36228 44402
rect 36176 44338 36228 44344
rect 36372 44334 36400 44900
rect 36452 44804 36504 44810
rect 36452 44746 36504 44752
rect 35716 44328 35768 44334
rect 35716 44270 35768 44276
rect 36360 44328 36412 44334
rect 36360 44270 36412 44276
rect 35532 43716 35584 43722
rect 35532 43658 35584 43664
rect 36464 43314 36492 44746
rect 36740 43382 36768 45426
rect 37200 45422 37228 45750
rect 37278 45656 37334 45665
rect 37278 45591 37334 45600
rect 37188 45416 37240 45422
rect 37188 45358 37240 45364
rect 37188 44736 37240 44742
rect 37188 44678 37240 44684
rect 36728 43376 36780 43382
rect 36728 43318 36780 43324
rect 36452 43308 36504 43314
rect 36452 43250 36504 43256
rect 34612 42764 34664 42770
rect 34612 42706 34664 42712
rect 34704 42764 34756 42770
rect 34704 42706 34756 42712
rect 35440 42764 35492 42770
rect 35440 42706 35492 42712
rect 34336 42696 34388 42702
rect 34336 42638 34388 42644
rect 34348 42362 34376 42638
rect 33968 42356 34020 42362
rect 33968 42298 34020 42304
rect 34336 42356 34388 42362
rect 34336 42298 34388 42304
rect 33980 41818 34008 42298
rect 36740 42294 36768 43318
rect 37200 42702 37228 44678
rect 37292 43994 37320 45591
rect 37384 45554 37412 46378
rect 37556 46028 37608 46034
rect 37556 45970 37608 45976
rect 37384 45526 37504 45554
rect 37372 45348 37424 45354
rect 37372 45290 37424 45296
rect 37384 44878 37412 45290
rect 37372 44872 37424 44878
rect 37372 44814 37424 44820
rect 37280 43988 37332 43994
rect 37280 43930 37332 43936
rect 37476 43382 37504 45526
rect 37568 45354 37596 45970
rect 37660 45966 37688 47058
rect 37844 46918 37872 49200
rect 37832 46912 37884 46918
rect 37832 46854 37884 46860
rect 38212 46714 38240 49200
rect 38476 47184 38528 47190
rect 38476 47126 38528 47132
rect 38384 47048 38436 47054
rect 38384 46990 38436 46996
rect 38200 46708 38252 46714
rect 38200 46650 38252 46656
rect 38396 46510 38424 46990
rect 38488 46578 38516 47126
rect 38580 47036 38608 49200
rect 38660 47048 38712 47054
rect 38580 47008 38660 47036
rect 38476 46572 38528 46578
rect 38476 46514 38528 46520
rect 38108 46504 38160 46510
rect 38108 46446 38160 46452
rect 38384 46504 38436 46510
rect 38384 46446 38436 46452
rect 37648 45960 37700 45966
rect 37648 45902 37700 45908
rect 38120 45898 38148 46446
rect 38488 46034 38516 46514
rect 38476 46028 38528 46034
rect 38476 45970 38528 45976
rect 38580 45966 38608 47008
rect 38660 46990 38712 46996
rect 38948 46374 38976 49200
rect 38936 46368 38988 46374
rect 38936 46310 38988 46316
rect 39316 46170 39344 49200
rect 39408 46986 39436 49286
rect 39670 49200 39726 49286
rect 40038 49314 40094 50000
rect 40038 49286 40356 49314
rect 40038 49200 40094 49286
rect 40224 47048 40276 47054
rect 40224 46990 40276 46996
rect 39396 46980 39448 46986
rect 39396 46922 39448 46928
rect 39948 46912 40000 46918
rect 39948 46854 40000 46860
rect 39580 46572 39632 46578
rect 39580 46514 39632 46520
rect 39488 46504 39540 46510
rect 39488 46446 39540 46452
rect 39304 46164 39356 46170
rect 39304 46106 39356 46112
rect 39500 46034 39528 46446
rect 39488 46028 39540 46034
rect 39488 45970 39540 45976
rect 38568 45960 38620 45966
rect 38568 45902 38620 45908
rect 39120 45960 39172 45966
rect 39120 45902 39172 45908
rect 38108 45892 38160 45898
rect 38108 45834 38160 45840
rect 38200 45892 38252 45898
rect 38200 45834 38252 45840
rect 38120 45490 38148 45834
rect 38108 45484 38160 45490
rect 38108 45426 38160 45432
rect 37648 45416 37700 45422
rect 37648 45358 37700 45364
rect 37556 45348 37608 45354
rect 37556 45290 37608 45296
rect 37660 45286 37688 45358
rect 37648 45280 37700 45286
rect 37648 45222 37700 45228
rect 37556 44872 37608 44878
rect 37660 44860 37688 45222
rect 37608 44832 37688 44860
rect 37556 44814 37608 44820
rect 37464 43376 37516 43382
rect 37464 43318 37516 43324
rect 37568 42770 37596 44814
rect 38120 43858 38148 45426
rect 38212 45422 38240 45834
rect 39132 45490 39160 45902
rect 38660 45484 38712 45490
rect 38660 45426 38712 45432
rect 39120 45484 39172 45490
rect 39120 45426 39172 45432
rect 38200 45416 38252 45422
rect 38200 45358 38252 45364
rect 38568 45416 38620 45422
rect 38568 45358 38620 45364
rect 38292 45348 38344 45354
rect 38292 45290 38344 45296
rect 38304 44402 38332 45290
rect 38292 44396 38344 44402
rect 38292 44338 38344 44344
rect 38476 44328 38528 44334
rect 38476 44270 38528 44276
rect 38488 43994 38516 44270
rect 38476 43988 38528 43994
rect 38476 43930 38528 43936
rect 38108 43852 38160 43858
rect 38108 43794 38160 43800
rect 37556 42764 37608 42770
rect 37556 42706 37608 42712
rect 37188 42696 37240 42702
rect 37188 42638 37240 42644
rect 36912 42560 36964 42566
rect 36912 42502 36964 42508
rect 36924 42362 36952 42502
rect 36912 42356 36964 42362
rect 36912 42298 36964 42304
rect 36728 42288 36780 42294
rect 36728 42230 36780 42236
rect 37200 42022 37228 42638
rect 38120 42362 38148 43794
rect 38580 43790 38608 45358
rect 38672 44878 38700 45426
rect 39304 45280 39356 45286
rect 39304 45222 39356 45228
rect 39316 44878 39344 45222
rect 39500 44946 39528 45970
rect 39592 45966 39620 46514
rect 39580 45960 39632 45966
rect 39580 45902 39632 45908
rect 39856 45348 39908 45354
rect 39856 45290 39908 45296
rect 39488 44940 39540 44946
rect 39488 44882 39540 44888
rect 38660 44872 38712 44878
rect 38660 44814 38712 44820
rect 39304 44872 39356 44878
rect 39304 44814 39356 44820
rect 38672 43790 38700 44814
rect 39868 44538 39896 45290
rect 39960 45082 39988 46854
rect 40236 46578 40264 46990
rect 40328 46578 40356 49286
rect 40406 49200 40462 50000
rect 40774 49314 40830 50000
rect 40512 49286 40830 49314
rect 40420 47258 40448 49200
rect 40408 47252 40460 47258
rect 40408 47194 40460 47200
rect 40224 46572 40276 46578
rect 40224 46514 40276 46520
rect 40316 46572 40368 46578
rect 40316 46514 40368 46520
rect 40132 45892 40184 45898
rect 40132 45834 40184 45840
rect 39948 45076 40000 45082
rect 39948 45018 40000 45024
rect 39856 44532 39908 44538
rect 39856 44474 39908 44480
rect 39948 44328 40000 44334
rect 39948 44270 40000 44276
rect 39396 44192 39448 44198
rect 39396 44134 39448 44140
rect 38568 43784 38620 43790
rect 38568 43726 38620 43732
rect 38660 43784 38712 43790
rect 38660 43726 38712 43732
rect 39408 43314 39436 44134
rect 39960 43314 39988 44270
rect 39396 43308 39448 43314
rect 39396 43250 39448 43256
rect 39948 43308 40000 43314
rect 39948 43250 40000 43256
rect 40144 42770 40172 45834
rect 40512 45554 40540 49286
rect 40774 49200 40830 49286
rect 41142 49200 41198 50000
rect 41510 49200 41566 50000
rect 41878 49200 41934 50000
rect 42246 49314 42302 50000
rect 42246 49286 42564 49314
rect 42246 49200 42302 49286
rect 40592 46912 40644 46918
rect 40592 46854 40644 46860
rect 40604 46034 40632 46854
rect 40684 46504 40736 46510
rect 40682 46472 40684 46481
rect 40736 46472 40738 46481
rect 40682 46407 40738 46416
rect 41156 46102 41184 49200
rect 41420 46708 41472 46714
rect 41420 46650 41472 46656
rect 41432 46322 41460 46650
rect 41524 46510 41552 49200
rect 41788 47184 41840 47190
rect 41788 47126 41840 47132
rect 41512 46504 41564 46510
rect 41512 46446 41564 46452
rect 41432 46294 41552 46322
rect 41144 46096 41196 46102
rect 41144 46038 41196 46044
rect 40592 46028 40644 46034
rect 40592 45970 40644 45976
rect 40776 45960 40828 45966
rect 40776 45902 40828 45908
rect 41236 45960 41288 45966
rect 41236 45902 41288 45908
rect 40592 45620 40644 45626
rect 40592 45562 40644 45568
rect 40236 45526 40540 45554
rect 40236 44742 40264 45526
rect 40316 45484 40368 45490
rect 40316 45426 40368 45432
rect 40328 44946 40356 45426
rect 40604 45422 40632 45562
rect 40788 45490 40816 45902
rect 41248 45626 41276 45902
rect 41420 45824 41472 45830
rect 41420 45766 41472 45772
rect 41236 45620 41288 45626
rect 41236 45562 41288 45568
rect 40776 45484 40828 45490
rect 40776 45426 40828 45432
rect 40408 45416 40460 45422
rect 40408 45358 40460 45364
rect 40592 45416 40644 45422
rect 40592 45358 40644 45364
rect 40316 44940 40368 44946
rect 40316 44882 40368 44888
rect 40224 44736 40276 44742
rect 40224 44678 40276 44684
rect 40420 44470 40448 45358
rect 40408 44464 40460 44470
rect 40408 44406 40460 44412
rect 40604 44402 40632 45358
rect 40788 44810 40816 45426
rect 41248 44860 41276 45562
rect 41432 44946 41460 45766
rect 41524 45490 41552 46294
rect 41800 45558 41828 47126
rect 41788 45552 41840 45558
rect 41788 45494 41840 45500
rect 41512 45484 41564 45490
rect 41512 45426 41564 45432
rect 41420 44940 41472 44946
rect 41420 44882 41472 44888
rect 41328 44872 41380 44878
rect 41248 44832 41328 44860
rect 41328 44814 41380 44820
rect 40776 44804 40828 44810
rect 40776 44746 40828 44752
rect 40788 44402 40816 44746
rect 41340 44538 41368 44814
rect 41328 44532 41380 44538
rect 41328 44474 41380 44480
rect 40592 44396 40644 44402
rect 40592 44338 40644 44344
rect 40776 44396 40828 44402
rect 40776 44338 40828 44344
rect 40604 43994 40632 44338
rect 41892 44266 41920 49200
rect 42432 47048 42484 47054
rect 42432 46990 42484 46996
rect 42444 46889 42472 46990
rect 42430 46880 42486 46889
rect 42430 46815 42486 46824
rect 42248 46028 42300 46034
rect 42248 45970 42300 45976
rect 42260 45898 42288 45970
rect 42248 45892 42300 45898
rect 42248 45834 42300 45840
rect 42260 45082 42288 45834
rect 42536 45554 42564 49286
rect 42614 49200 42670 50000
rect 42982 49200 43038 50000
rect 43350 49200 43406 50000
rect 43718 49314 43774 50000
rect 43718 49286 44036 49314
rect 43718 49200 43774 49286
rect 42628 46170 42656 49200
rect 42616 46164 42668 46170
rect 42616 46106 42668 46112
rect 42996 46073 43024 49200
rect 43260 47048 43312 47054
rect 43260 46990 43312 46996
rect 43272 46753 43300 46990
rect 43258 46744 43314 46753
rect 43258 46679 43314 46688
rect 43364 46578 43392 49200
rect 44008 47274 44036 49286
rect 44086 49200 44142 50000
rect 44454 49314 44510 50000
rect 44454 49286 44772 49314
rect 44454 49200 44510 49286
rect 44100 47410 44128 49200
rect 44100 47382 44312 47410
rect 44008 47258 44220 47274
rect 44008 47252 44232 47258
rect 44008 47246 44180 47252
rect 44180 47194 44232 47200
rect 44284 47190 44312 47382
rect 44272 47184 44324 47190
rect 44272 47126 44324 47132
rect 43904 46912 43956 46918
rect 43904 46854 43956 46860
rect 43352 46572 43404 46578
rect 43352 46514 43404 46520
rect 42982 46064 43038 46073
rect 42982 45999 43038 46008
rect 43916 45626 43944 46854
rect 44284 46170 44312 47126
rect 44744 46918 44772 49286
rect 44822 49200 44878 50000
rect 45190 49200 45246 50000
rect 45558 49314 45614 50000
rect 45558 49286 45876 49314
rect 45558 49200 45614 49286
rect 44732 46912 44784 46918
rect 44732 46854 44784 46860
rect 44836 46578 44864 49200
rect 44824 46572 44876 46578
rect 44824 46514 44876 46520
rect 44272 46164 44324 46170
rect 44272 46106 44324 46112
rect 45204 45626 45232 49200
rect 45848 46578 45876 49286
rect 45926 49200 45982 50000
rect 45940 47258 45968 49200
rect 45928 47252 45980 47258
rect 45928 47194 45980 47200
rect 45836 46572 45888 46578
rect 45836 46514 45888 46520
rect 43904 45620 43956 45626
rect 43904 45562 43956 45568
rect 45192 45620 45244 45626
rect 45192 45562 45244 45568
rect 42536 45526 42656 45554
rect 42628 45490 42656 45526
rect 42616 45484 42668 45490
rect 42616 45426 42668 45432
rect 43260 45416 43312 45422
rect 43260 45358 43312 45364
rect 42708 45280 42760 45286
rect 42708 45222 42760 45228
rect 42248 45076 42300 45082
rect 42248 45018 42300 45024
rect 42260 44538 42288 45018
rect 42720 44946 42748 45222
rect 42708 44940 42760 44946
rect 42708 44882 42760 44888
rect 43272 44742 43300 45358
rect 43260 44736 43312 44742
rect 43260 44678 43312 44684
rect 42248 44532 42300 44538
rect 42248 44474 42300 44480
rect 41880 44260 41932 44266
rect 41880 44202 41932 44208
rect 43272 43994 43300 44678
rect 40592 43988 40644 43994
rect 40592 43930 40644 43936
rect 43260 43988 43312 43994
rect 43260 43930 43312 43936
rect 41144 43648 41196 43654
rect 41144 43590 41196 43596
rect 41156 42770 41184 43590
rect 40132 42764 40184 42770
rect 40132 42706 40184 42712
rect 41144 42764 41196 42770
rect 41144 42706 41196 42712
rect 38108 42356 38160 42362
rect 38108 42298 38160 42304
rect 35532 42016 35584 42022
rect 35532 41958 35584 41964
rect 37188 42016 37240 42022
rect 37188 41958 37240 41964
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 33968 41812 34020 41818
rect 33968 41754 34020 41760
rect 35544 41750 35572 41958
rect 33140 41744 33192 41750
rect 33140 41686 33192 41692
rect 35532 41744 35584 41750
rect 35532 41686 35584 41692
rect 32404 41268 32456 41274
rect 32404 41210 32456 41216
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 31024 3664 31076 3670
rect 31024 3606 31076 3612
rect 30840 3460 30892 3466
rect 30840 3402 30892 3408
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 30760 800 30788 2382
rect 31036 800 31064 3606
rect 31852 3528 31904 3534
rect 31852 3470 31904 3476
rect 32680 3528 32732 3534
rect 32680 3470 32732 3476
rect 33232 3528 33284 3534
rect 33232 3470 33284 3476
rect 35348 3528 35400 3534
rect 35348 3470 35400 3476
rect 35440 3528 35492 3534
rect 35440 3470 35492 3476
rect 36268 3528 36320 3534
rect 36268 3470 36320 3476
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 37924 3528 37976 3534
rect 37924 3470 37976 3476
rect 39028 3528 39080 3534
rect 39028 3470 39080 3476
rect 40408 3528 40460 3534
rect 40408 3470 40460 3476
rect 40960 3528 41012 3534
rect 40960 3470 41012 3476
rect 41512 3528 41564 3534
rect 41512 3470 41564 3476
rect 42892 3528 42944 3534
rect 42892 3470 42944 3476
rect 43168 3528 43220 3534
rect 43168 3470 43220 3476
rect 44824 3528 44876 3534
rect 44824 3470 44876 3476
rect 45652 3528 45704 3534
rect 45652 3470 45704 3476
rect 46480 3528 46532 3534
rect 46480 3470 46532 3476
rect 46756 3528 46808 3534
rect 46756 3470 46808 3476
rect 47308 3528 47360 3534
rect 47308 3470 47360 3476
rect 31208 2984 31260 2990
rect 31208 2926 31260 2932
rect 31220 2650 31248 2926
rect 31300 2848 31352 2854
rect 31300 2790 31352 2796
rect 31208 2644 31260 2650
rect 31208 2586 31260 2592
rect 31312 800 31340 2790
rect 31576 2508 31628 2514
rect 31576 2450 31628 2456
rect 31588 800 31616 2450
rect 31864 800 31892 3470
rect 32404 2848 32456 2854
rect 32404 2790 32456 2796
rect 32128 2576 32180 2582
rect 32128 2518 32180 2524
rect 32140 800 32168 2518
rect 32416 800 32444 2790
rect 32692 800 32720 3470
rect 32956 2984 33008 2990
rect 32956 2926 33008 2932
rect 32968 800 32996 2926
rect 33244 800 33272 3470
rect 34796 2916 34848 2922
rect 34796 2858 34848 2864
rect 33784 2848 33836 2854
rect 33784 2790 33836 2796
rect 34336 2848 34388 2854
rect 34336 2790 34388 2796
rect 33508 2508 33560 2514
rect 33508 2450 33560 2456
rect 33520 800 33548 2450
rect 33796 800 33824 2790
rect 34060 2440 34112 2446
rect 34060 2382 34112 2388
rect 34072 800 34100 2382
rect 34348 800 34376 2790
rect 34612 2576 34664 2582
rect 34612 2518 34664 2524
rect 34624 800 34652 2518
rect 34808 1442 34836 2858
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 1850 35388 3470
rect 35176 1822 35388 1850
rect 34808 1414 34928 1442
rect 34900 800 34928 1414
rect 35176 800 35204 1822
rect 35452 800 35480 3470
rect 35716 2848 35768 2854
rect 35716 2790 35768 2796
rect 35728 800 35756 2790
rect 35992 2440 36044 2446
rect 35992 2382 36044 2388
rect 36004 800 36032 2382
rect 36280 800 36308 3470
rect 36820 2848 36872 2854
rect 36820 2790 36872 2796
rect 36544 2508 36596 2514
rect 36544 2450 36596 2456
rect 36556 800 36584 2450
rect 36832 800 36860 2790
rect 37108 800 37136 3470
rect 37648 2848 37700 2854
rect 37648 2790 37700 2796
rect 37372 2372 37424 2378
rect 37372 2314 37424 2320
rect 37384 800 37412 2314
rect 37660 800 37688 2790
rect 37936 800 37964 3470
rect 38752 2984 38804 2990
rect 38752 2926 38804 2932
rect 38200 2848 38252 2854
rect 38200 2790 38252 2796
rect 38212 800 38240 2790
rect 38476 2576 38528 2582
rect 38476 2518 38528 2524
rect 38488 800 38516 2518
rect 38764 800 38792 2926
rect 39040 800 39068 3470
rect 39580 2848 39632 2854
rect 39580 2790 39632 2796
rect 40132 2848 40184 2854
rect 40132 2790 40184 2796
rect 39304 2508 39356 2514
rect 39304 2450 39356 2456
rect 39316 800 39344 2450
rect 39592 800 39620 2790
rect 39856 2440 39908 2446
rect 39856 2382 39908 2388
rect 39868 800 39896 2382
rect 40144 800 40172 2790
rect 40420 800 40448 3470
rect 40684 2984 40736 2990
rect 40684 2926 40736 2932
rect 40696 800 40724 2926
rect 40972 800 41000 3470
rect 41236 2508 41288 2514
rect 41236 2450 41288 2456
rect 41248 800 41276 2450
rect 41524 800 41552 3470
rect 42616 2984 42668 2990
rect 42616 2926 42668 2932
rect 42064 2848 42116 2854
rect 42064 2790 42116 2796
rect 41788 2440 41840 2446
rect 41788 2382 41840 2388
rect 41800 800 41828 2382
rect 42076 800 42104 2790
rect 42340 2576 42392 2582
rect 42340 2518 42392 2524
rect 42352 800 42380 2518
rect 42628 800 42656 2926
rect 42904 800 42932 3470
rect 43180 800 43208 3470
rect 44548 2984 44600 2990
rect 44548 2926 44600 2932
rect 43444 2848 43496 2854
rect 43444 2790 43496 2796
rect 43996 2848 44048 2854
rect 43996 2790 44048 2796
rect 43456 800 43484 2790
rect 43720 2508 43772 2514
rect 43720 2450 43772 2456
rect 43732 800 43760 2450
rect 44008 800 44036 2790
rect 44272 2372 44324 2378
rect 44272 2314 44324 2320
rect 44284 800 44312 2314
rect 44560 800 44588 2926
rect 44836 800 44864 3470
rect 45376 2848 45428 2854
rect 45376 2790 45428 2796
rect 45100 2576 45152 2582
rect 45100 2518 45152 2524
rect 45112 800 45140 2518
rect 45388 800 45416 2790
rect 45664 800 45692 3470
rect 45928 2848 45980 2854
rect 45928 2790 45980 2796
rect 45940 800 45968 2790
rect 46204 2440 46256 2446
rect 46204 2382 46256 2388
rect 46216 800 46244 2382
rect 46492 800 46520 3470
rect 46768 800 46796 3470
rect 47032 2848 47084 2854
rect 47032 2790 47084 2796
rect 47044 800 47072 2790
rect 47320 800 47348 3470
rect 2410 0 2466 800
rect 2502 0 2558 800
rect 2594 0 2650 800
rect 2686 0 2742 800
rect 2778 0 2834 800
rect 2870 0 2926 800
rect 2962 0 3018 800
rect 3054 0 3110 800
rect 3146 0 3202 800
rect 3238 0 3294 800
rect 3330 0 3386 800
rect 3422 0 3478 800
rect 3514 0 3570 800
rect 3606 0 3662 800
rect 3698 0 3754 800
rect 3790 0 3846 800
rect 3882 0 3938 800
rect 3974 0 4030 800
rect 4066 0 4122 800
rect 4158 0 4214 800
rect 4250 0 4306 800
rect 4342 0 4398 800
rect 4434 0 4490 800
rect 4526 0 4582 800
rect 4618 0 4674 800
rect 4710 0 4766 800
rect 4802 0 4858 800
rect 4894 0 4950 800
rect 4986 0 5042 800
rect 5078 0 5134 800
rect 5170 0 5226 800
rect 5262 0 5318 800
rect 5354 0 5410 800
rect 5446 0 5502 800
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5722 0 5778 800
rect 5814 0 5870 800
rect 5906 0 5962 800
rect 5998 0 6054 800
rect 6090 0 6146 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6366 0 6422 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6642 0 6698 800
rect 6734 0 6790 800
rect 6826 0 6882 800
rect 6918 0 6974 800
rect 7010 0 7066 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7286 0 7342 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
<< via2 >>
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 18970 46572 19026 46608
rect 18970 46552 18972 46572
rect 18972 46552 19024 46572
rect 19024 46552 19026 46572
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19338 46436 19394 46472
rect 19338 46416 19340 46436
rect 19340 46416 19392 46436
rect 19392 46416 19394 46436
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 20902 46280 20958 46336
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 21822 46688 21878 46744
rect 22098 46688 22154 46744
rect 22834 46416 22890 46472
rect 22098 46280 22154 46336
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 29550 46008 29606 46064
rect 30470 46824 30526 46880
rect 33598 46688 33654 46744
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34334 46416 34390 46472
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 35530 46572 35586 46608
rect 35530 46552 35532 46572
rect 35532 46552 35584 46572
rect 35584 46552 35586 46572
rect 36358 46824 36414 46880
rect 36726 46824 36782 46880
rect 37186 46688 37242 46744
rect 37094 45600 37150 45656
rect 37278 45600 37334 45656
rect 40682 46452 40684 46472
rect 40684 46452 40736 46472
rect 40736 46452 40738 46472
rect 40682 46416 40738 46452
rect 42430 46824 42486 46880
rect 43258 46688 43314 46744
rect 42982 46008 43038 46064
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
<< metal3 >>
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 30465 46882 30531 46885
rect 36353 46882 36419 46885
rect 30465 46880 36419 46882
rect 30465 46824 30470 46880
rect 30526 46824 36358 46880
rect 36414 46824 36419 46880
rect 30465 46822 36419 46824
rect 30465 46819 30531 46822
rect 36353 46819 36419 46822
rect 36721 46882 36787 46885
rect 42425 46882 42491 46885
rect 36721 46880 42491 46882
rect 36721 46824 36726 46880
rect 36782 46824 42430 46880
rect 42486 46824 42491 46880
rect 36721 46822 42491 46824
rect 36721 46819 36787 46822
rect 42425 46819 42491 46822
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 21817 46746 21883 46749
rect 22093 46746 22159 46749
rect 33593 46746 33659 46749
rect 21817 46744 33659 46746
rect 21817 46688 21822 46744
rect 21878 46688 22098 46744
rect 22154 46688 33598 46744
rect 33654 46688 33659 46744
rect 21817 46686 33659 46688
rect 21817 46683 21883 46686
rect 22093 46683 22159 46686
rect 33593 46683 33659 46686
rect 37181 46746 37247 46749
rect 43253 46746 43319 46749
rect 37181 46744 43319 46746
rect 37181 46688 37186 46744
rect 37242 46688 43258 46744
rect 43314 46688 43319 46744
rect 37181 46686 43319 46688
rect 37181 46683 37247 46686
rect 43253 46683 43319 46686
rect 18965 46610 19031 46613
rect 35525 46610 35591 46613
rect 18965 46608 35591 46610
rect 18965 46552 18970 46608
rect 19026 46552 35530 46608
rect 35586 46552 35591 46608
rect 18965 46550 35591 46552
rect 18965 46547 19031 46550
rect 35525 46547 35591 46550
rect 19333 46474 19399 46477
rect 22829 46474 22895 46477
rect 19333 46472 22895 46474
rect 19333 46416 19338 46472
rect 19394 46416 22834 46472
rect 22890 46416 22895 46472
rect 19333 46414 22895 46416
rect 19333 46411 19399 46414
rect 22829 46411 22895 46414
rect 34329 46474 34395 46477
rect 40677 46474 40743 46477
rect 34329 46472 40743 46474
rect 34329 46416 34334 46472
rect 34390 46416 40682 46472
rect 40738 46416 40743 46472
rect 34329 46414 40743 46416
rect 34329 46411 34395 46414
rect 40677 46411 40743 46414
rect 20897 46338 20963 46341
rect 22093 46338 22159 46341
rect 20897 46336 22159 46338
rect 20897 46280 20902 46336
rect 20958 46280 22098 46336
rect 22154 46280 22159 46336
rect 20897 46278 22159 46280
rect 20897 46275 20963 46278
rect 22093 46275 22159 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 29545 46066 29611 46069
rect 42977 46066 43043 46069
rect 29545 46064 43043 46066
rect 29545 46008 29550 46064
rect 29606 46008 42982 46064
rect 43038 46008 43043 46064
rect 29545 46006 43043 46008
rect 29545 46003 29611 46006
rect 42977 46003 43043 46006
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 37089 45658 37155 45661
rect 37273 45658 37339 45661
rect 37089 45656 37339 45658
rect 37089 45600 37094 45656
rect 37150 45600 37278 45656
rect 37334 45600 37339 45656
rect 37089 45598 37339 45600
rect 37089 45595 37155 45598
rect 37273 45595 37339 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 20148 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A
timestamp 1666199351
transform 1 0 21252 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A
timestamp 1666199351
transform -1 0 19596 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A
timestamp 1666199351
transform -1 0 32476 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A_N
timestamp 1666199351
transform 1 0 31280 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__B
timestamp 1666199351
transform 1 0 32292 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A1
timestamp 1666199351
transform -1 0 31280 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A2
timestamp 1666199351
transform -1 0 31556 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A
timestamp 1666199351
transform 1 0 26496 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A
timestamp 1666199351
transform -1 0 20700 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A1
timestamp 1666199351
transform 1 0 31188 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1666199351
transform -1 0 30176 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 1666199351
transform 1 0 26128 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A
timestamp 1666199351
transform -1 0 28888 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A1
timestamp 1666199351
transform 1 0 29624 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__B1_N
timestamp 1666199351
transform -1 0 31832 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__B1
timestamp 1666199351
transform -1 0 27876 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A
timestamp 1666199351
transform -1 0 35144 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A
timestamp 1666199351
transform -1 0 31924 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 1666199351
transform 1 0 22632 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A
timestamp 1666199351
transform 1 0 25944 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A1
timestamp 1666199351
transform 1 0 30544 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A
timestamp 1666199351
transform -1 0 20148 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A
timestamp 1666199351
transform -1 0 39284 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A_N
timestamp 1666199351
transform 1 0 43792 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__B
timestamp 1666199351
transform 1 0 44252 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A1
timestamp 1666199351
transform -1 0 37628 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A2
timestamp 1666199351
transform -1 0 36524 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1666199351
transform -1 0 35052 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1666199351
transform -1 0 34316 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A1
timestamp 1666199351
transform -1 0 38180 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A
timestamp 1666199351
transform 1 0 37444 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1666199351
transform -1 0 35144 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A
timestamp 1666199351
transform -1 0 41492 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A1
timestamp 1666199351
transform -1 0 38732 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__B1_N
timestamp 1666199351
transform -1 0 41308 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__B1
timestamp 1666199351
transform -1 0 40204 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A
timestamp 1666199351
transform -1 0 40756 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1666199351
transform 1 0 39284 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A
timestamp 1666199351
transform 1 0 33764 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A
timestamp 1666199351
transform -1 0 34592 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A1
timestamp 1666199351
transform 1 0 37444 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A
timestamp 1666199351
transform 1 0 43240 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1666199351
transform 1 0 27876 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A2_N
timestamp 1666199351
transform 1 0 29716 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__B2
timestamp 1666199351
transform 1 0 33396 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A2
timestamp 1666199351
transform -1 0 26680 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A3
timestamp 1666199351
transform -1 0 26128 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A
timestamp 1666199351
transform -1 0 41860 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A2_N
timestamp 1666199351
transform 1 0 42688 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__B2
timestamp 1666199351
transform -1 0 42780 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A2
timestamp 1666199351
transform 1 0 41860 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A3
timestamp 1666199351
transform -1 0 43424 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__B
timestamp 1666199351
transform -1 0 16376 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A
timestamp 1666199351
transform -1 0 17296 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__A2_N
timestamp 1666199351
transform -1 0 18400 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A
timestamp 1666199351
transform -1 0 29256 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A2
timestamp 1666199351
transform -1 0 25024 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__B1
timestamp 1666199351
transform -1 0 25576 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A
timestamp 1666199351
transform -1 0 44712 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__A2
timestamp 1666199351
transform 1 0 42136 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__B1
timestamp 1666199351
transform -1 0 38180 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A2
timestamp 1666199351
transform -1 0 27324 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__B1
timestamp 1666199351
transform 1 0 27140 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__B
timestamp 1666199351
transform -1 0 24472 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A
timestamp 1666199351
transform -1 0 28244 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__B1
timestamp 1666199351
transform 1 0 30820 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A1
timestamp 1666199351
transform -1 0 28704 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__A2
timestamp 1666199351
transform -1 0 36248 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__B1
timestamp 1666199351
transform -1 0 36800 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__B
timestamp 1666199351
transform -1 0 33396 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A
timestamp 1666199351
transform -1 0 37076 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__A1
timestamp 1666199351
transform -1 0 25208 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__B1
timestamp 1666199351
transform -1 0 25024 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A1
timestamp 1666199351
transform -1 0 19596 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A1
timestamp 1666199351
transform 1 0 35512 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__B1
timestamp 1666199351
transform -1 0 42136 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__A1
timestamp 1666199351
transform 1 0 33120 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__C1
timestamp 1666199351
transform 1 0 19596 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19
timestamp 1666199351
transform 1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40
timestamp 1666199351
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47
timestamp 1666199351
transform 1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1666199351
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1666199351
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1666199351
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1666199351
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1666199351
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1666199351
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1666199351
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1666199351
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1666199351
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1666199351
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124
timestamp 1666199351
transform 1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131
timestamp 1666199351
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1666199351
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1666199351
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152
timestamp 1666199351
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_159
timestamp 1666199351
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1666199351
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1666199351
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_180
timestamp 1666199351
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1666199351
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1666199351
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1666199351
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1666199351
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1666199351
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1666199351
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1666199351
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1666199351
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1666199351
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1666199351
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_257
timestamp 1666199351
transform 1 0 24748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_271
timestamp 1666199351
transform 1 0 26036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1666199351
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_281
timestamp 1666199351
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_287
timestamp 1666199351
transform 1 0 27508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1666199351
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1666199351
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1666199351
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_316
timestamp 1666199351
transform 1 0 30176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_323
timestamp 1666199351
transform 1 0 30820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1666199351
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1666199351
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_342
timestamp 1666199351
transform 1 0 32568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1666199351
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1666199351
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1666199351
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_370
timestamp 1666199351
transform 1 0 35144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1666199351
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1666199351
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1666199351
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_398
timestamp 1666199351
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_405
timestamp 1666199351
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 1666199351
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1666199351
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_426
timestamp 1666199351
transform 1 0 40296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_433
timestamp 1666199351
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_440
timestamp 1666199351
transform 1 0 41584 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1666199351
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_454
timestamp 1666199351
transform 1 0 42872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 1666199351
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_468
timestamp 1666199351
transform 1 0 44160 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1666199351
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_482
timestamp 1666199351
transform 1 0 45448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_489
timestamp 1666199351
transform 1 0 46092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_496
timestamp 1666199351
transform 1 0 46736 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1666199351
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_510
timestamp 1666199351
transform 1 0 48024 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_15
timestamp 1666199351
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_19
timestamp 1666199351
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp 1666199351
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_33
timestamp 1666199351
transform 1 0 4140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1666199351
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_47
timestamp 1666199351
transform 1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1666199351
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1666199351
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_68
timestamp 1666199351
transform 1 0 7360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_75
timestamp 1666199351
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1666199351
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_89
timestamp 1666199351
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1666199351
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1666199351
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1666199351
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1666199351
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_124
timestamp 1666199351
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_131
timestamp 1666199351
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_138
timestamp 1666199351
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1666199351
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_152
timestamp 1666199351
transform 1 0 15088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_159
timestamp 1666199351
transform 1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1666199351
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_169
timestamp 1666199351
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1666199351
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1666199351
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_194
timestamp 1666199351
transform 1 0 18952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_201
timestamp 1666199351
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_210
timestamp 1666199351
transform 1 0 20424 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_216
timestamp 1666199351
transform 1 0 20976 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1666199351
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1666199351
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_240
timestamp 1666199351
transform 1 0 23184 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_244
timestamp 1666199351
transform 1 0 23552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_258
timestamp 1666199351
transform 1 0 24840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_275
timestamp 1666199351
transform 1 0 26404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1666199351
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1666199351
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_296
timestamp 1666199351
transform 1 0 28336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_313
timestamp 1666199351
transform 1 0 29900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_322
timestamp 1666199351
transform 1 0 30728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1666199351
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1666199351
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1666199351
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_342
timestamp 1666199351
transform 1 0 32568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_349
timestamp 1666199351
transform 1 0 33212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_356
timestamp 1666199351
transform 1 0 33856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_363
timestamp 1666199351
transform 1 0 34500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_370
timestamp 1666199351
transform 1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_377
timestamp 1666199351
transform 1 0 35788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_384
timestamp 1666199351
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1666199351
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_398
timestamp 1666199351
transform 1 0 37720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_405
timestamp 1666199351
transform 1 0 38364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_412
timestamp 1666199351
transform 1 0 39008 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_419
timestamp 1666199351
transform 1 0 39652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_426
timestamp 1666199351
transform 1 0 40296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_433
timestamp 1666199351
transform 1 0 40940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_440
timestamp 1666199351
transform 1 0 41584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1666199351
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_454
timestamp 1666199351
transform 1 0 42872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1666199351
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_468
timestamp 1666199351
transform 1 0 44160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_475
timestamp 1666199351
transform 1 0 44804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_482
timestamp 1666199351
transform 1 0 45448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_489
timestamp 1666199351
transform 1 0 46092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_496
timestamp 1666199351
transform 1 0 46736 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1666199351
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_510
timestamp 1666199351
transform 1 0 48024 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666199351
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666199351
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666199351
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_35
timestamp 1666199351
transform 1 0 4324 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1666199351
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_45
timestamp 1666199351
transform 1 0 5244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_54
timestamp 1666199351
transform 1 0 6072 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_63
timestamp 1666199351
transform 1 0 6900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_72
timestamp 1666199351
transform 1 0 7728 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1666199351
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1666199351
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_90
timestamp 1666199351
transform 1 0 9384 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_99
timestamp 1666199351
transform 1 0 10212 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1666199351
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_112
timestamp 1666199351
transform 1 0 11408 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_116
timestamp 1666199351
transform 1 0 11776 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_123
timestamp 1666199351
transform 1 0 12420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_130
timestamp 1666199351
transform 1 0 13064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1666199351
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1666199351
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_152
timestamp 1666199351
transform 1 0 15088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1666199351
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_166
timestamp 1666199351
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1666199351
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1666199351
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_187
timestamp 1666199351
transform 1 0 18308 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1666199351
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1666199351
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_201
timestamp 1666199351
transform 1 0 19596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_218
timestamp 1666199351
transform 1 0 21160 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_227
timestamp 1666199351
transform 1 0 21988 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_244
timestamp 1666199351
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_253
timestamp 1666199351
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_266
timestamp 1666199351
transform 1 0 25576 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_274
timestamp 1666199351
transform 1 0 26312 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_280
timestamp 1666199351
transform 1 0 26864 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_288
timestamp 1666199351
transform 1 0 27600 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp 1666199351
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1666199351
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1666199351
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_314
timestamp 1666199351
transform 1 0 29992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1666199351
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_328
timestamp 1666199351
transform 1 0 31280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_335
timestamp 1666199351
transform 1 0 31924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_342
timestamp 1666199351
transform 1 0 32568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_349
timestamp 1666199351
transform 1 0 33212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_356
timestamp 1666199351
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_365
timestamp 1666199351
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_371
timestamp 1666199351
transform 1 0 35236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_378
timestamp 1666199351
transform 1 0 35880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_385
timestamp 1666199351
transform 1 0 36524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_392
timestamp 1666199351
transform 1 0 37168 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_401
timestamp 1666199351
transform 1 0 37996 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_409
timestamp 1666199351
transform 1 0 38732 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1666199351
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1666199351
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_421
timestamp 1666199351
transform 1 0 39836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_428
timestamp 1666199351
transform 1 0 40480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_435
timestamp 1666199351
transform 1 0 41124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_442
timestamp 1666199351
transform 1 0 41768 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_450
timestamp 1666199351
transform 1 0 42504 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_455
timestamp 1666199351
transform 1 0 42964 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_462
timestamp 1666199351
transform 1 0 43608 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 1666199351
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1666199351
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_482
timestamp 1666199351
transform 1 0 45448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_489
timestamp 1666199351
transform 1 0 46092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_496
timestamp 1666199351
transform 1 0 46736 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_503
timestamp 1666199351
transform 1 0 47380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_510
timestamp 1666199351
transform 1 0 48024 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666199351
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666199351
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666199351
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666199351
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1666199351
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666199351
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666199351
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666199351
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666199351
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666199351
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666199351
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666199351
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666199351
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666199351
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666199351
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666199351
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1666199351
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1666199351
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_176
timestamp 1666199351
transform 1 0 17296 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_183
timestamp 1666199351
transform 1 0 17940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_190
timestamp 1666199351
transform 1 0 18584 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_197
timestamp 1666199351
transform 1 0 19228 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_204
timestamp 1666199351
transform 1 0 19872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_213
timestamp 1666199351
transform 1 0 20700 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1666199351
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1666199351
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_240
timestamp 1666199351
transform 1 0 23184 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_257
timestamp 1666199351
transform 1 0 24748 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_268
timestamp 1666199351
transform 1 0 25760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_272
timestamp 1666199351
transform 1 0 26128 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1666199351
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1666199351
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_296
timestamp 1666199351
transform 1 0 28336 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_305
timestamp 1666199351
transform 1 0 29164 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_312
timestamp 1666199351
transform 1 0 29808 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_319
timestamp 1666199351
transform 1 0 30452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_331
timestamp 1666199351
transform 1 0 31556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1666199351
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1666199351
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1666199351
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1666199351
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1666199351
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1666199351
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1666199351
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1666199351
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1666199351
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1666199351
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1666199351
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1666199351
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1666199351
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1666199351
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1666199351
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1666199351
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1666199351
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1666199351
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1666199351
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_505
timestamp 1666199351
transform 1 0 47564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_513
timestamp 1666199351
transform 1 0 48300 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666199351
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666199351
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666199351
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666199351
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666199351
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666199351
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666199351
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666199351
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666199351
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666199351
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666199351
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666199351
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666199351
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666199351
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666199351
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666199351
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666199351
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666199351
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_177
timestamp 1666199351
transform 1 0 17388 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_183
timestamp 1666199351
transform 1 0 17940 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_187
timestamp 1666199351
transform 1 0 18308 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1666199351
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1666199351
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_204
timestamp 1666199351
transform 1 0 19872 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_213
timestamp 1666199351
transform 1 0 20700 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_230
timestamp 1666199351
transform 1 0 22264 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_241
timestamp 1666199351
transform 1 0 23276 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1666199351
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1666199351
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_258
timestamp 1666199351
transform 1 0 24840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_275
timestamp 1666199351
transform 1 0 26404 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_283
timestamp 1666199351
transform 1 0 27140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_287
timestamp 1666199351
transform 1 0 27508 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1666199351
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1666199351
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_316
timestamp 1666199351
transform 1 0 30176 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_323
timestamp 1666199351
transform 1 0 30820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_335
timestamp 1666199351
transform 1 0 31924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_347
timestamp 1666199351
transform 1 0 33028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_359
timestamp 1666199351
transform 1 0 34132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1666199351
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1666199351
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1666199351
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1666199351
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1666199351
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1666199351
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1666199351
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1666199351
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1666199351
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1666199351
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1666199351
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1666199351
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1666199351
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1666199351
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1666199351
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1666199351
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_513
timestamp 1666199351
transform 1 0 48300 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666199351
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666199351
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1666199351
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1666199351
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1666199351
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666199351
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666199351
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666199351
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666199351
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666199351
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666199351
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666199351
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666199351
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666199351
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666199351
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666199351
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666199351
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666199351
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666199351
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666199351
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1666199351
transform 1 0 18860 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_198
timestamp 1666199351
transform 1 0 19320 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1666199351
transform 1 0 20884 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1666199351
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_225
timestamp 1666199351
transform 1 0 21804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_231
timestamp 1666199351
transform 1 0 22356 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_245
timestamp 1666199351
transform 1 0 23644 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_249
timestamp 1666199351
transform 1 0 24012 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_263
timestamp 1666199351
transform 1 0 25300 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_271
timestamp 1666199351
transform 1 0 26036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1666199351
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1666199351
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_296
timestamp 1666199351
transform 1 0 28336 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_313
timestamp 1666199351
transform 1 0 29900 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_325
timestamp 1666199351
transform 1 0 31004 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_333
timestamp 1666199351
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1666199351
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1666199351
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1666199351
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1666199351
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1666199351
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1666199351
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1666199351
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1666199351
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1666199351
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1666199351
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1666199351
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1666199351
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1666199351
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1666199351
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1666199351
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1666199351
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1666199351
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1666199351
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_505
timestamp 1666199351
transform 1 0 47564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_513
timestamp 1666199351
transform 1 0 48300 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666199351
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666199351
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666199351
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666199351
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666199351
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666199351
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666199351
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666199351
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666199351
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666199351
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666199351
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666199351
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666199351
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666199351
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666199351
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666199351
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666199351
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666199351
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666199351
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666199351
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666199351
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_197
timestamp 1666199351
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_208
timestamp 1666199351
transform 1 0 20240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_212
timestamp 1666199351
transform 1 0 20608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_218
timestamp 1666199351
transform 1 0 21160 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_222
timestamp 1666199351
transform 1 0 21528 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_228
timestamp 1666199351
transform 1 0 22080 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_237
timestamp 1666199351
transform 1 0 22908 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1666199351
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1666199351
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_260
timestamp 1666199351
transform 1 0 25024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_269
timestamp 1666199351
transform 1 0 25852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_277
timestamp 1666199351
transform 1 0 26588 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_283
timestamp 1666199351
transform 1 0 27140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_297
timestamp 1666199351
transform 1 0 28428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1666199351
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1666199351
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1666199351
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1666199351
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1666199351
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1666199351
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1666199351
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1666199351
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1666199351
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1666199351
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1666199351
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1666199351
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1666199351
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1666199351
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1666199351
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1666199351
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1666199351
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1666199351
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1666199351
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1666199351
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1666199351
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1666199351
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_513
timestamp 1666199351
transform 1 0 48300 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666199351
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666199351
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666199351
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1666199351
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1666199351
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666199351
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666199351
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666199351
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666199351
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666199351
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666199351
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666199351
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666199351
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666199351
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666199351
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666199351
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666199351
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666199351
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666199351
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666199351
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_193
timestamp 1666199351
transform 1 0 18860 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_201
timestamp 1666199351
transform 1 0 19596 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_205
timestamp 1666199351
transform 1 0 19964 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1666199351
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1666199351
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 1666199351
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_261
timestamp 1666199351
transform 1 0 25116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1666199351
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_281
timestamp 1666199351
transform 1 0 26956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_290
timestamp 1666199351
transform 1 0 27784 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_299
timestamp 1666199351
transform 1 0 28612 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_306
timestamp 1666199351
transform 1 0 29256 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_318
timestamp 1666199351
transform 1 0 30360 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_330
timestamp 1666199351
transform 1 0 31464 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1666199351
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1666199351
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1666199351
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1666199351
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1666199351
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1666199351
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1666199351
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1666199351
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1666199351
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1666199351
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1666199351
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1666199351
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1666199351
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1666199351
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1666199351
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1666199351
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1666199351
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1666199351
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_505
timestamp 1666199351
transform 1 0 47564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_513
timestamp 1666199351
transform 1 0 48300 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666199351
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666199351
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666199351
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666199351
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666199351
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666199351
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666199351
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666199351
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666199351
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666199351
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666199351
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666199351
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666199351
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666199351
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666199351
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666199351
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666199351
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666199351
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666199351
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666199351
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666199351
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1666199351
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_205
timestamp 1666199351
transform 1 0 19964 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1666199351
transform 1 0 20332 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_217
timestamp 1666199351
transform 1 0 21068 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_225
timestamp 1666199351
transform 1 0 21804 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_233
timestamp 1666199351
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1666199351
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1666199351
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_260
timestamp 1666199351
transform 1 0 25024 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_271
timestamp 1666199351
transform 1 0 26036 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_279
timestamp 1666199351
transform 1 0 26772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_287
timestamp 1666199351
transform 1 0 27508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1666199351
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1666199351
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1666199351
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1666199351
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1666199351
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1666199351
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1666199351
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1666199351
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1666199351
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1666199351
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1666199351
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1666199351
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1666199351
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1666199351
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1666199351
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1666199351
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1666199351
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1666199351
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1666199351
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1666199351
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1666199351
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1666199351
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1666199351
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_513
timestamp 1666199351
transform 1 0 48300 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666199351
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666199351
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1666199351
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1666199351
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1666199351
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666199351
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666199351
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666199351
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666199351
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666199351
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666199351
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666199351
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666199351
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666199351
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666199351
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666199351
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666199351
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666199351
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666199351
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666199351
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666199351
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666199351
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_217
timestamp 1666199351
transform 1 0 21068 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1666199351
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1666199351
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_230
timestamp 1666199351
transform 1 0 22264 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_239
timestamp 1666199351
transform 1 0 23092 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_247
timestamp 1666199351
transform 1 0 23828 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_261
timestamp 1666199351
transform 1 0 25116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1666199351
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1666199351
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_286
timestamp 1666199351
transform 1 0 27416 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1666199351
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1666199351
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1666199351
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1666199351
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1666199351
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1666199351
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1666199351
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1666199351
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1666199351
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1666199351
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1666199351
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1666199351
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1666199351
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1666199351
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1666199351
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1666199351
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1666199351
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1666199351
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1666199351
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1666199351
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1666199351
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1666199351
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1666199351
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_505
timestamp 1666199351
transform 1 0 47564 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_513
timestamp 1666199351
transform 1 0 48300 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666199351
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666199351
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666199351
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666199351
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666199351
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666199351
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666199351
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666199351
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666199351
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666199351
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666199351
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666199351
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666199351
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666199351
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666199351
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666199351
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666199351
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666199351
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666199351
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666199351
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666199351
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666199351
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666199351
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666199351
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_233
timestamp 1666199351
transform 1 0 22540 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_238
timestamp 1666199351
transform 1 0 23000 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_246
timestamp 1666199351
transform 1 0 23736 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1666199351
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1666199351
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_258
timestamp 1666199351
transform 1 0 24840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_262
timestamp 1666199351
transform 1 0 25208 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_267
timestamp 1666199351
transform 1 0 25668 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_274
timestamp 1666199351
transform 1 0 26312 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_286
timestamp 1666199351
transform 1 0 27416 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_298
timestamp 1666199351
transform 1 0 28520 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1666199351
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1666199351
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1666199351
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1666199351
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1666199351
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1666199351
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1666199351
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1666199351
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1666199351
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1666199351
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1666199351
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1666199351
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1666199351
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1666199351
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1666199351
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1666199351
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1666199351
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1666199351
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1666199351
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1666199351
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1666199351
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1666199351
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_513
timestamp 1666199351
transform 1 0 48300 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666199351
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666199351
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666199351
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666199351
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666199351
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666199351
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666199351
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666199351
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666199351
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666199351
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666199351
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666199351
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666199351
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666199351
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666199351
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666199351
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666199351
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666199351
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666199351
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666199351
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666199351
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666199351
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666199351
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666199351
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1666199351
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1666199351
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1666199351
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1666199351
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1666199351
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1666199351
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666199351
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1666199351
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1666199351
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1666199351
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1666199351
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1666199351
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1666199351
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1666199351
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1666199351
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1666199351
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1666199351
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1666199351
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1666199351
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1666199351
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1666199351
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1666199351
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1666199351
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1666199351
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1666199351
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1666199351
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1666199351
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1666199351
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1666199351
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1666199351
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1666199351
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1666199351
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666199351
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666199351
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666199351
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666199351
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666199351
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666199351
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666199351
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666199351
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666199351
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666199351
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666199351
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666199351
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666199351
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666199351
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666199351
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666199351
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666199351
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666199351
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666199351
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666199351
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666199351
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666199351
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666199351
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1666199351
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1666199351
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1666199351
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1666199351
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1666199351
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1666199351
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1666199351
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1666199351
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1666199351
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1666199351
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1666199351
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1666199351
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1666199351
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1666199351
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1666199351
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1666199351
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1666199351
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1666199351
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1666199351
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1666199351
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1666199351
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1666199351
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1666199351
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1666199351
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1666199351
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1666199351
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1666199351
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1666199351
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1666199351
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1666199351
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1666199351
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_513
timestamp 1666199351
transform 1 0 48300 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666199351
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1666199351
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1666199351
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1666199351
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1666199351
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1666199351
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666199351
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666199351
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666199351
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666199351
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666199351
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666199351
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666199351
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666199351
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666199351
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666199351
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666199351
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666199351
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666199351
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666199351
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666199351
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1666199351
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1666199351
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666199351
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666199351
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666199351
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666199351
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666199351
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1666199351
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666199351
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1666199351
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1666199351
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1666199351
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1666199351
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1666199351
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1666199351
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1666199351
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1666199351
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1666199351
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1666199351
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1666199351
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1666199351
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1666199351
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1666199351
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1666199351
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1666199351
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1666199351
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1666199351
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1666199351
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1666199351
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1666199351
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1666199351
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1666199351
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1666199351
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1666199351
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1666199351
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1666199351
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1666199351
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666199351
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666199351
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666199351
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666199351
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666199351
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666199351
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666199351
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666199351
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666199351
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666199351
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666199351
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666199351
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666199351
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666199351
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666199351
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666199351
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666199351
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666199351
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666199351
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666199351
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1666199351
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1666199351
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1666199351
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1666199351
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1666199351
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1666199351
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1666199351
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1666199351
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1666199351
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1666199351
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1666199351
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1666199351
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1666199351
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1666199351
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1666199351
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1666199351
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1666199351
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1666199351
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1666199351
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1666199351
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1666199351
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1666199351
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1666199351
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1666199351
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1666199351
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1666199351
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1666199351
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1666199351
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1666199351
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1666199351
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1666199351
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1666199351
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_513
timestamp 1666199351
transform 1 0 48300 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666199351
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666199351
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666199351
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1666199351
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1666199351
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666199351
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666199351
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666199351
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666199351
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666199351
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666199351
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666199351
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666199351
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666199351
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666199351
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666199351
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666199351
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666199351
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666199351
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666199351
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666199351
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666199351
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666199351
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666199351
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666199351
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1666199351
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1666199351
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666199351
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1666199351
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666199351
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1666199351
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1666199351
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1666199351
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1666199351
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1666199351
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1666199351
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1666199351
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1666199351
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1666199351
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1666199351
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1666199351
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1666199351
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1666199351
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1666199351
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1666199351
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1666199351
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1666199351
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1666199351
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1666199351
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1666199351
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1666199351
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1666199351
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1666199351
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1666199351
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_505
timestamp 1666199351
transform 1 0 47564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_513
timestamp 1666199351
transform 1 0 48300 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666199351
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666199351
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666199351
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666199351
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666199351
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666199351
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666199351
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666199351
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666199351
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666199351
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666199351
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666199351
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666199351
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666199351
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666199351
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666199351
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666199351
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666199351
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666199351
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1666199351
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666199351
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666199351
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666199351
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666199351
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1666199351
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1666199351
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666199351
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666199351
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1666199351
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1666199351
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1666199351
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1666199351
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1666199351
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1666199351
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1666199351
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1666199351
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1666199351
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1666199351
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1666199351
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1666199351
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1666199351
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1666199351
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1666199351
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1666199351
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1666199351
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1666199351
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1666199351
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1666199351
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1666199351
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1666199351
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1666199351
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1666199351
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1666199351
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1666199351
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_513
timestamp 1666199351
transform 1 0 48300 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1666199351
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666199351
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1666199351
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1666199351
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1666199351
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1666199351
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666199351
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666199351
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666199351
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666199351
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666199351
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666199351
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666199351
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666199351
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666199351
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666199351
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666199351
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666199351
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666199351
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666199351
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666199351
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666199351
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666199351
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666199351
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1666199351
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1666199351
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1666199351
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1666199351
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1666199351
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666199351
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1666199351
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1666199351
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1666199351
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1666199351
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1666199351
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1666199351
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1666199351
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1666199351
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1666199351
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1666199351
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1666199351
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1666199351
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1666199351
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1666199351
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1666199351
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1666199351
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1666199351
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1666199351
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1666199351
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1666199351
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1666199351
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1666199351
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1666199351
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1666199351
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1666199351
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_513
timestamp 1666199351
transform 1 0 48300 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666199351
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1666199351
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666199351
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666199351
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666199351
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666199351
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666199351
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666199351
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666199351
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666199351
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666199351
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666199351
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666199351
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666199351
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666199351
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666199351
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666199351
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1666199351
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1666199351
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1666199351
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666199351
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666199351
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666199351
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1666199351
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1666199351
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1666199351
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666199351
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1666199351
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1666199351
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1666199351
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1666199351
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1666199351
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1666199351
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1666199351
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1666199351
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1666199351
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1666199351
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1666199351
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1666199351
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1666199351
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1666199351
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1666199351
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1666199351
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1666199351
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1666199351
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1666199351
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1666199351
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1666199351
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1666199351
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1666199351
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1666199351
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1666199351
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1666199351
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1666199351
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1666199351
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666199351
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666199351
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666199351
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666199351
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1666199351
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666199351
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666199351
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666199351
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666199351
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666199351
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666199351
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666199351
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666199351
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666199351
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666199351
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666199351
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1666199351
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666199351
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666199351
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666199351
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666199351
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666199351
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666199351
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666199351
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666199351
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1666199351
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1666199351
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1666199351
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1666199351
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1666199351
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1666199351
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1666199351
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1666199351
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1666199351
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1666199351
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1666199351
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1666199351
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1666199351
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1666199351
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1666199351
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1666199351
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1666199351
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1666199351
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1666199351
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1666199351
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1666199351
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1666199351
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1666199351
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1666199351
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1666199351
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1666199351
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1666199351
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1666199351
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1666199351
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1666199351
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1666199351
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1666199351
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1666199351
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666199351
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666199351
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666199351
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666199351
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666199351
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666199351
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666199351
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666199351
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666199351
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666199351
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666199351
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666199351
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666199351
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666199351
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666199351
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1666199351
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1666199351
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1666199351
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666199351
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666199351
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666199351
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1666199351
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1666199351
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1666199351
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1666199351
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1666199351
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1666199351
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1666199351
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1666199351
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1666199351
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1666199351
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1666199351
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1666199351
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1666199351
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1666199351
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1666199351
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1666199351
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1666199351
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1666199351
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1666199351
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1666199351
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1666199351
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1666199351
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1666199351
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1666199351
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1666199351
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1666199351
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1666199351
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1666199351
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1666199351
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1666199351
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1666199351
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_513
timestamp 1666199351
transform 1 0 48300 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666199351
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666199351
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666199351
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666199351
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666199351
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666199351
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666199351
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666199351
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666199351
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666199351
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666199351
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666199351
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666199351
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666199351
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666199351
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666199351
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666199351
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666199351
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666199351
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666199351
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666199351
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1666199351
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666199351
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666199351
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1666199351
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1666199351
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1666199351
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1666199351
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1666199351
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666199351
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1666199351
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1666199351
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1666199351
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1666199351
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1666199351
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1666199351
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1666199351
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1666199351
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1666199351
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1666199351
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1666199351
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1666199351
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1666199351
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1666199351
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1666199351
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1666199351
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1666199351
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1666199351
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1666199351
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1666199351
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1666199351
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1666199351
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1666199351
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1666199351
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1666199351
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_513
timestamp 1666199351
transform 1 0 48300 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666199351
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1666199351
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666199351
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666199351
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666199351
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666199351
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666199351
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666199351
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666199351
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666199351
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666199351
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666199351
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666199351
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666199351
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666199351
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666199351
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666199351
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666199351
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666199351
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666199351
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666199351
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666199351
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666199351
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1666199351
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1666199351
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1666199351
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1666199351
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1666199351
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1666199351
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1666199351
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1666199351
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1666199351
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1666199351
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1666199351
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1666199351
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1666199351
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1666199351
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1666199351
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1666199351
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1666199351
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1666199351
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1666199351
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1666199351
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1666199351
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1666199351
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1666199351
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1666199351
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1666199351
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1666199351
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1666199351
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1666199351
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1666199351
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1666199351
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1666199351
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1666199351
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666199351
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666199351
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666199351
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1666199351
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1666199351
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666199351
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666199351
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666199351
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666199351
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666199351
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666199351
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666199351
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666199351
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666199351
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666199351
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666199351
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666199351
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666199351
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666199351
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666199351
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666199351
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666199351
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666199351
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666199351
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1666199351
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1666199351
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1666199351
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1666199351
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1666199351
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1666199351
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1666199351
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1666199351
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1666199351
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1666199351
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1666199351
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1666199351
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1666199351
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1666199351
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1666199351
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1666199351
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1666199351
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1666199351
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1666199351
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1666199351
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1666199351
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1666199351
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1666199351
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1666199351
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1666199351
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1666199351
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1666199351
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1666199351
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1666199351
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1666199351
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1666199351
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1666199351
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666199351
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1666199351
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666199351
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666199351
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666199351
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666199351
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666199351
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666199351
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666199351
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666199351
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666199351
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666199351
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666199351
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666199351
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666199351
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666199351
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666199351
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666199351
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666199351
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666199351
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666199351
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666199351
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666199351
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1666199351
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1666199351
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1666199351
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1666199351
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1666199351
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1666199351
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1666199351
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1666199351
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1666199351
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1666199351
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1666199351
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1666199351
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1666199351
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1666199351
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1666199351
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1666199351
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1666199351
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1666199351
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1666199351
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1666199351
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1666199351
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1666199351
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1666199351
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1666199351
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1666199351
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1666199351
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1666199351
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1666199351
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1666199351
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1666199351
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1666199351
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_513
timestamp 1666199351
transform 1 0 48300 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666199351
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666199351
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666199351
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1666199351
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1666199351
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666199351
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666199351
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666199351
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666199351
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666199351
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666199351
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666199351
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666199351
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666199351
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666199351
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666199351
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666199351
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666199351
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666199351
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666199351
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666199351
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666199351
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666199351
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666199351
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1666199351
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1666199351
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1666199351
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1666199351
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1666199351
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1666199351
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1666199351
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1666199351
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1666199351
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1666199351
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1666199351
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1666199351
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1666199351
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1666199351
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1666199351
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1666199351
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1666199351
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1666199351
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1666199351
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1666199351
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1666199351
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1666199351
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1666199351
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1666199351
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1666199351
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1666199351
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1666199351
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1666199351
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1666199351
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1666199351
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_505
timestamp 1666199351
transform 1 0 47564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_513
timestamp 1666199351
transform 1 0 48300 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666199351
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666199351
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666199351
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666199351
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666199351
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666199351
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666199351
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666199351
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666199351
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666199351
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666199351
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666199351
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666199351
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666199351
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666199351
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666199351
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666199351
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666199351
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666199351
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666199351
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666199351
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666199351
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666199351
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1666199351
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1666199351
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1666199351
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1666199351
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1666199351
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1666199351
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1666199351
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1666199351
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1666199351
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1666199351
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1666199351
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1666199351
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1666199351
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1666199351
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1666199351
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1666199351
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1666199351
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1666199351
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1666199351
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1666199351
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1666199351
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1666199351
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1666199351
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1666199351
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1666199351
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1666199351
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1666199351
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1666199351
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1666199351
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1666199351
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1666199351
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_513
timestamp 1666199351
transform 1 0 48300 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666199351
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666199351
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666199351
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666199351
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1666199351
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666199351
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666199351
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666199351
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666199351
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666199351
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666199351
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666199351
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666199351
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666199351
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666199351
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666199351
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666199351
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666199351
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666199351
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666199351
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666199351
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666199351
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666199351
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666199351
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1666199351
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1666199351
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1666199351
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1666199351
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1666199351
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1666199351
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1666199351
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1666199351
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1666199351
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1666199351
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1666199351
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1666199351
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1666199351
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1666199351
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1666199351
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1666199351
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1666199351
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1666199351
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1666199351
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1666199351
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1666199351
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1666199351
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1666199351
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1666199351
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1666199351
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1666199351
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1666199351
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1666199351
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1666199351
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1666199351
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1666199351
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_513
timestamp 1666199351
transform 1 0 48300 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666199351
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1666199351
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666199351
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666199351
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666199351
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666199351
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666199351
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666199351
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666199351
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666199351
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666199351
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666199351
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666199351
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666199351
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666199351
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666199351
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666199351
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666199351
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666199351
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666199351
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666199351
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666199351
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666199351
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1666199351
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1666199351
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1666199351
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1666199351
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1666199351
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1666199351
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1666199351
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1666199351
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1666199351
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1666199351
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1666199351
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1666199351
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1666199351
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1666199351
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1666199351
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1666199351
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1666199351
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1666199351
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1666199351
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1666199351
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1666199351
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1666199351
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1666199351
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1666199351
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1666199351
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1666199351
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1666199351
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1666199351
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1666199351
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1666199351
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1666199351
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_513
timestamp 1666199351
transform 1 0 48300 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1666199351
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1666199351
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1666199351
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1666199351
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1666199351
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1666199351
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666199351
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666199351
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666199351
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666199351
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666199351
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666199351
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666199351
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666199351
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666199351
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666199351
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666199351
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666199351
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666199351
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666199351
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666199351
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666199351
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666199351
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666199351
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1666199351
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1666199351
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1666199351
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1666199351
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1666199351
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1666199351
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1666199351
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1666199351
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1666199351
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1666199351
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1666199351
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1666199351
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1666199351
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1666199351
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1666199351
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1666199351
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1666199351
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1666199351
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1666199351
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1666199351
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1666199351
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1666199351
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1666199351
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1666199351
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1666199351
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1666199351
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1666199351
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1666199351
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1666199351
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1666199351
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1666199351
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_513
timestamp 1666199351
transform 1 0 48300 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666199351
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666199351
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666199351
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666199351
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666199351
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666199351
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666199351
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666199351
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666199351
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666199351
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666199351
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666199351
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666199351
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666199351
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666199351
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666199351
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666199351
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666199351
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1666199351
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666199351
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666199351
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666199351
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666199351
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1666199351
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1666199351
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1666199351
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1666199351
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1666199351
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1666199351
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1666199351
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1666199351
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1666199351
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1666199351
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1666199351
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1666199351
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1666199351
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1666199351
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1666199351
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1666199351
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1666199351
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1666199351
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1666199351
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1666199351
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1666199351
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1666199351
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1666199351
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1666199351
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1666199351
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1666199351
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1666199351
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1666199351
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1666199351
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1666199351
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1666199351
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_513
timestamp 1666199351
transform 1 0 48300 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666199351
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666199351
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666199351
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666199351
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1666199351
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666199351
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666199351
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666199351
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666199351
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666199351
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666199351
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666199351
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666199351
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666199351
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666199351
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666199351
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666199351
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666199351
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666199351
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666199351
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666199351
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666199351
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1666199351
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666199351
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1666199351
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1666199351
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1666199351
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1666199351
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1666199351
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1666199351
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1666199351
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1666199351
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1666199351
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1666199351
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1666199351
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1666199351
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1666199351
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1666199351
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1666199351
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1666199351
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1666199351
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1666199351
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1666199351
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1666199351
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1666199351
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1666199351
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1666199351
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1666199351
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1666199351
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1666199351
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1666199351
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1666199351
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1666199351
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1666199351
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_505
timestamp 1666199351
transform 1 0 47564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_513
timestamp 1666199351
transform 1 0 48300 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666199351
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1666199351
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666199351
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666199351
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666199351
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666199351
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666199351
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666199351
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666199351
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666199351
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666199351
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666199351
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666199351
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666199351
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666199351
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666199351
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666199351
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666199351
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666199351
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1666199351
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666199351
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666199351
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1666199351
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1666199351
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1666199351
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1666199351
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1666199351
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1666199351
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1666199351
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1666199351
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1666199351
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1666199351
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1666199351
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1666199351
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1666199351
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1666199351
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1666199351
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1666199351
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1666199351
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1666199351
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1666199351
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1666199351
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1666199351
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1666199351
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1666199351
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1666199351
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1666199351
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1666199351
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1666199351
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1666199351
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1666199351
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1666199351
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1666199351
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1666199351
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_513
timestamp 1666199351
transform 1 0 48300 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666199351
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666199351
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1666199351
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1666199351
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1666199351
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666199351
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666199351
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666199351
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666199351
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666199351
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666199351
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666199351
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666199351
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666199351
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666199351
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666199351
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666199351
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666199351
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666199351
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666199351
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1666199351
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1666199351
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1666199351
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666199351
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1666199351
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1666199351
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1666199351
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1666199351
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1666199351
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1666199351
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1666199351
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1666199351
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1666199351
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1666199351
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1666199351
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1666199351
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1666199351
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1666199351
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1666199351
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1666199351
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1666199351
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1666199351
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1666199351
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1666199351
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1666199351
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1666199351
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1666199351
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1666199351
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1666199351
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1666199351
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1666199351
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1666199351
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1666199351
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1666199351
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1666199351
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_513
timestamp 1666199351
transform 1 0 48300 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666199351
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666199351
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666199351
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666199351
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666199351
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666199351
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666199351
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666199351
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666199351
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666199351
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666199351
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666199351
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666199351
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666199351
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666199351
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666199351
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666199351
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666199351
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666199351
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666199351
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666199351
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666199351
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1666199351
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1666199351
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1666199351
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1666199351
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1666199351
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1666199351
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1666199351
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1666199351
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1666199351
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1666199351
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1666199351
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1666199351
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1666199351
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1666199351
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1666199351
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1666199351
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1666199351
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1666199351
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1666199351
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1666199351
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1666199351
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1666199351
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1666199351
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1666199351
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1666199351
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1666199351
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1666199351
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1666199351
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1666199351
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1666199351
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1666199351
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1666199351
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_513
timestamp 1666199351
transform 1 0 48300 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666199351
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1666199351
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1666199351
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1666199351
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1666199351
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1666199351
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666199351
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666199351
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666199351
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666199351
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666199351
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666199351
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666199351
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666199351
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1666199351
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1666199351
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1666199351
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666199351
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666199351
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666199351
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1666199351
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1666199351
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1666199351
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1666199351
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1666199351
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1666199351
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1666199351
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1666199351
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1666199351
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1666199351
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1666199351
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1666199351
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1666199351
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1666199351
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1666199351
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1666199351
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1666199351
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1666199351
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1666199351
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1666199351
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1666199351
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1666199351
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1666199351
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1666199351
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1666199351
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1666199351
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1666199351
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1666199351
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1666199351
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1666199351
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1666199351
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1666199351
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1666199351
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1666199351
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1666199351
transform 1 0 47564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_513
timestamp 1666199351
transform 1 0 48300 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666199351
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666199351
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666199351
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666199351
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666199351
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666199351
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666199351
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666199351
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666199351
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666199351
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666199351
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666199351
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1666199351
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1666199351
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666199351
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666199351
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666199351
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666199351
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1666199351
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1666199351
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1666199351
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1666199351
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1666199351
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1666199351
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1666199351
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1666199351
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1666199351
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1666199351
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1666199351
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1666199351
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1666199351
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1666199351
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1666199351
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1666199351
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1666199351
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1666199351
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1666199351
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1666199351
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1666199351
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1666199351
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1666199351
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1666199351
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1666199351
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1666199351
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1666199351
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1666199351
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1666199351
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1666199351
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1666199351
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1666199351
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1666199351
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1666199351
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1666199351
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1666199351
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_513
timestamp 1666199351
transform 1 0 48300 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666199351
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1666199351
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1666199351
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1666199351
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1666199351
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1666199351
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666199351
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666199351
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666199351
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666199351
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666199351
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666199351
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666199351
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666199351
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666199351
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666199351
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666199351
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666199351
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1666199351
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1666199351
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1666199351
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1666199351
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1666199351
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666199351
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1666199351
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1666199351
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1666199351
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1666199351
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1666199351
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666199351
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1666199351
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1666199351
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1666199351
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1666199351
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1666199351
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1666199351
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1666199351
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1666199351
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1666199351
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1666199351
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1666199351
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1666199351
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1666199351
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1666199351
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1666199351
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1666199351
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1666199351
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1666199351
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1666199351
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1666199351
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1666199351
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1666199351
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1666199351
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1666199351
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1666199351
transform 1 0 47564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_513
timestamp 1666199351
transform 1 0 48300 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666199351
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1666199351
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666199351
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666199351
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666199351
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666199351
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666199351
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666199351
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666199351
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666199351
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666199351
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666199351
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666199351
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666199351
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666199351
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666199351
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1666199351
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1666199351
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1666199351
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1666199351
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666199351
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1666199351
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1666199351
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1666199351
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1666199351
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1666199351
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1666199351
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1666199351
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1666199351
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1666199351
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1666199351
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1666199351
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1666199351
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1666199351
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1666199351
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1666199351
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1666199351
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1666199351
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1666199351
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1666199351
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1666199351
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1666199351
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1666199351
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1666199351
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1666199351
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1666199351
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1666199351
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1666199351
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1666199351
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1666199351
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1666199351
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1666199351
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1666199351
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1666199351
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_513
timestamp 1666199351
transform 1 0 48300 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1666199351
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1666199351
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1666199351
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1666199351
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1666199351
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1666199351
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666199351
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666199351
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666199351
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666199351
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666199351
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666199351
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666199351
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666199351
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666199351
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1666199351
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1666199351
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666199351
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666199351
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1666199351
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1666199351
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1666199351
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1666199351
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666199351
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1666199351
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1666199351
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1666199351
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1666199351
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1666199351
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1666199351
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1666199351
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1666199351
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1666199351
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1666199351
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1666199351
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1666199351
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1666199351
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1666199351
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1666199351
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1666199351
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1666199351
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1666199351
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1666199351
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1666199351
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1666199351
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1666199351
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1666199351
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1666199351
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1666199351
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1666199351
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1666199351
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1666199351
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1666199351
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1666199351
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1666199351
transform 1 0 47564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_513
timestamp 1666199351
transform 1 0 48300 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1666199351
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1666199351
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666199351
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666199351
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666199351
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666199351
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666199351
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666199351
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666199351
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666199351
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666199351
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666199351
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666199351
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666199351
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666199351
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666199351
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1666199351
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1666199351
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1666199351
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1666199351
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1666199351
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666199351
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1666199351
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1666199351
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1666199351
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1666199351
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1666199351
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1666199351
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1666199351
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1666199351
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1666199351
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1666199351
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1666199351
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1666199351
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1666199351
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1666199351
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1666199351
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1666199351
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1666199351
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1666199351
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1666199351
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1666199351
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1666199351
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1666199351
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1666199351
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1666199351
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1666199351
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1666199351
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1666199351
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1666199351
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1666199351
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1666199351
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1666199351
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1666199351
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_513
timestamp 1666199351
transform 1 0 48300 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666199351
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666199351
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666199351
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666199351
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666199351
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666199351
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666199351
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1666199351
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1666199351
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1666199351
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1666199351
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666199351
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666199351
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1666199351
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1666199351
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1666199351
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1666199351
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1666199351
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666199351
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1666199351
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1666199351
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1666199351
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1666199351
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1666199351
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1666199351
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1666199351
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1666199351
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1666199351
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1666199351
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1666199351
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1666199351
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1666199351
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1666199351
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1666199351
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1666199351
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1666199351
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1666199351
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1666199351
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1666199351
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1666199351
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1666199351
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1666199351
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1666199351
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1666199351
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1666199351
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1666199351
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1666199351
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1666199351
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1666199351
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1666199351
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1666199351
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1666199351
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1666199351
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1666199351
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_505
timestamp 1666199351
transform 1 0 47564 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_513
timestamp 1666199351
transform 1 0 48300 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666199351
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1666199351
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666199351
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666199351
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1666199351
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1666199351
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666199351
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1666199351
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666199351
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666199351
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666199351
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1666199351
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1666199351
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1666199351
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666199351
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666199351
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1666199351
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1666199351
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1666199351
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1666199351
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1666199351
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1666199351
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1666199351
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1666199351
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1666199351
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1666199351
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666199351
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1666199351
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1666199351
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1666199351
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1666199351
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1666199351
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1666199351
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1666199351
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1666199351
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1666199351
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1666199351
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1666199351
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1666199351
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1666199351
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1666199351
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1666199351
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1666199351
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1666199351
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1666199351
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1666199351
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1666199351
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1666199351
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1666199351
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1666199351
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1666199351
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1666199351
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1666199351
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1666199351
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_513
timestamp 1666199351
transform 1 0 48300 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1666199351
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1666199351
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1666199351
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1666199351
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1666199351
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1666199351
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666199351
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666199351
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1666199351
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1666199351
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666199351
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666199351
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1666199351
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1666199351
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1666199351
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1666199351
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1666199351
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1666199351
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1666199351
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1666199351
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1666199351
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1666199351
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1666199351
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1666199351
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666199351
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1666199351
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1666199351
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1666199351
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1666199351
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1666199351
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1666199351
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1666199351
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1666199351
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1666199351
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1666199351
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1666199351
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1666199351
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1666199351
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1666199351
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1666199351
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1666199351
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1666199351
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1666199351
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1666199351
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1666199351
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1666199351
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1666199351
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1666199351
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1666199351
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1666199351
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1666199351
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1666199351
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1666199351
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1666199351
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_505
timestamp 1666199351
transform 1 0 47564 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_513
timestamp 1666199351
transform 1 0 48300 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1666199351
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1666199351
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666199351
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666199351
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666199351
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666199351
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666199351
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666199351
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666199351
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1666199351
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1666199351
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1666199351
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1666199351
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1666199351
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666199351
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666199351
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666199351
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1666199351
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1666199351
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1666199351
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1666199351
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1666199351
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1666199351
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1666199351
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1666199351
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1666199351
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666199351
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1666199351
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1666199351
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1666199351
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1666199351
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1666199351
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1666199351
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1666199351
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1666199351
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1666199351
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1666199351
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1666199351
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1666199351
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1666199351
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1666199351
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1666199351
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1666199351
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1666199351
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1666199351
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1666199351
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1666199351
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1666199351
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1666199351
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1666199351
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1666199351
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1666199351
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1666199351
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1666199351
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_513
timestamp 1666199351
transform 1 0 48300 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666199351
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666199351
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666199351
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666199351
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666199351
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666199351
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666199351
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666199351
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1666199351
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1666199351
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1666199351
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1666199351
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1666199351
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1666199351
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1666199351
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1666199351
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666199351
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666199351
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1666199351
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1666199351
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1666199351
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1666199351
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1666199351
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666199351
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1666199351
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1666199351
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1666199351
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1666199351
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1666199351
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1666199351
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1666199351
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1666199351
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1666199351
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1666199351
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1666199351
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1666199351
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1666199351
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1666199351
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1666199351
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1666199351
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1666199351
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1666199351
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1666199351
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1666199351
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1666199351
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1666199351
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1666199351
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1666199351
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1666199351
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1666199351
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1666199351
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1666199351
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1666199351
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1666199351
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1666199351
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1666199351
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666199351
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666199351
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666199351
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666199351
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666199351
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1666199351
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1666199351
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1666199351
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666199351
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1666199351
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1666199351
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1666199351
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1666199351
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1666199351
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666199351
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1666199351
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1666199351
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1666199351
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1666199351
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1666199351
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1666199351
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666199351
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1666199351
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1666199351
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1666199351
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1666199351
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1666199351
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1666199351
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1666199351
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1666199351
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1666199351
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1666199351
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1666199351
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1666199351
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1666199351
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1666199351
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1666199351
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1666199351
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1666199351
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1666199351
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1666199351
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1666199351
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1666199351
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1666199351
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1666199351
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1666199351
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1666199351
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1666199351
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1666199351
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1666199351
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1666199351
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1666199351
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1666199351
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1666199351
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_513
timestamp 1666199351
transform 1 0 48300 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666199351
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666199351
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666199351
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1666199351
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1666199351
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1666199351
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666199351
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1666199351
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1666199351
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1666199351
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1666199351
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1666199351
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1666199351
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1666199351
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1666199351
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1666199351
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1666199351
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1666199351
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1666199351
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1666199351
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1666199351
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1666199351
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1666199351
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1666199351
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1666199351
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1666199351
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1666199351
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1666199351
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1666199351
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1666199351
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1666199351
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1666199351
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1666199351
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1666199351
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1666199351
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1666199351
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1666199351
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1666199351
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1666199351
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1666199351
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1666199351
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1666199351
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1666199351
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1666199351
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1666199351
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1666199351
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1666199351
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1666199351
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1666199351
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1666199351
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1666199351
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1666199351
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1666199351
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1666199351
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_505
timestamp 1666199351
transform 1 0 47564 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_513
timestamp 1666199351
transform 1 0 48300 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666199351
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1666199351
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666199351
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666199351
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666199351
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666199351
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666199351
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1666199351
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666199351
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1666199351
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1666199351
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1666199351
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1666199351
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1666199351
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666199351
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1666199351
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1666199351
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1666199351
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1666199351
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1666199351
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1666199351
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1666199351
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1666199351
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1666199351
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1666199351
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1666199351
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1666199351
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1666199351
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1666199351
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1666199351
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1666199351
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1666199351
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1666199351
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1666199351
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1666199351
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1666199351
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1666199351
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1666199351
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1666199351
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1666199351
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1666199351
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1666199351
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1666199351
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1666199351
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1666199351
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1666199351
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1666199351
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1666199351
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1666199351
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1666199351
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1666199351
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1666199351
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1666199351
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1666199351
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_513
timestamp 1666199351
transform 1 0 48300 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666199351
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666199351
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666199351
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666199351
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1666199351
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666199351
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666199351
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1666199351
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1666199351
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1666199351
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1666199351
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1666199351
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1666199351
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1666199351
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1666199351
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1666199351
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1666199351
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666199351
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1666199351
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1666199351
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1666199351
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1666199351
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1666199351
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1666199351
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1666199351
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1666199351
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1666199351
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1666199351
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1666199351
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1666199351
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1666199351
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1666199351
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1666199351
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1666199351
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1666199351
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1666199351
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1666199351
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1666199351
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1666199351
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1666199351
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1666199351
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1666199351
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1666199351
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1666199351
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1666199351
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1666199351
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1666199351
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1666199351
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1666199351
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1666199351
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1666199351
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1666199351
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1666199351
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1666199351
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1666199351
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1666199351
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666199351
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666199351
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666199351
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666199351
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666199351
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666199351
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666199351
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666199351
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666199351
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1666199351
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1666199351
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1666199351
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1666199351
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1666199351
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1666199351
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1666199351
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1666199351
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1666199351
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1666199351
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1666199351
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1666199351
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1666199351
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1666199351
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1666199351
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1666199351
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1666199351
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1666199351
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1666199351
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1666199351
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1666199351
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1666199351
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1666199351
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1666199351
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1666199351
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1666199351
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1666199351
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1666199351
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1666199351
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1666199351
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1666199351
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1666199351
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1666199351
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1666199351
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1666199351
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1666199351
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1666199351
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1666199351
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1666199351
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1666199351
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1666199351
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1666199351
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1666199351
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1666199351
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1666199351
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_513
timestamp 1666199351
transform 1 0 48300 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666199351
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666199351
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666199351
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666199351
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666199351
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666199351
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666199351
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666199351
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666199351
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666199351
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1666199351
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666199351
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666199351
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1666199351
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1666199351
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1666199351
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1666199351
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1666199351
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1666199351
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1666199351
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1666199351
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1666199351
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1666199351
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1666199351
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1666199351
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1666199351
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1666199351
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1666199351
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1666199351
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1666199351
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1666199351
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1666199351
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1666199351
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1666199351
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1666199351
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1666199351
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1666199351
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1666199351
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1666199351
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1666199351
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1666199351
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1666199351
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1666199351
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1666199351
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1666199351
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1666199351
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1666199351
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1666199351
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1666199351
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1666199351
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1666199351
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1666199351
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1666199351
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1666199351
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1666199351
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1666199351
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666199351
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1666199351
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666199351
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666199351
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666199351
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666199351
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666199351
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666199351
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666199351
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1666199351
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1666199351
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1666199351
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1666199351
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1666199351
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1666199351
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1666199351
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1666199351
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1666199351
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1666199351
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1666199351
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1666199351
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1666199351
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1666199351
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1666199351
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1666199351
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1666199351
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1666199351
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1666199351
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1666199351
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1666199351
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1666199351
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1666199351
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1666199351
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1666199351
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1666199351
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1666199351
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1666199351
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1666199351
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1666199351
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1666199351
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1666199351
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1666199351
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1666199351
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1666199351
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1666199351
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1666199351
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1666199351
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1666199351
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1666199351
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1666199351
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1666199351
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1666199351
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1666199351
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1666199351
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1666199351
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1666199351
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666199351
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1666199351
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1666199351
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1666199351
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1666199351
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666199351
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666199351
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1666199351
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1666199351
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1666199351
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1666199351
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666199351
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1666199351
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1666199351
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1666199351
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1666199351
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1666199351
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1666199351
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1666199351
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1666199351
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1666199351
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1666199351
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1666199351
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1666199351
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1666199351
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1666199351
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1666199351
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1666199351
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1666199351
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1666199351
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1666199351
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1666199351
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1666199351
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1666199351
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1666199351
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1666199351
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1666199351
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1666199351
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1666199351
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1666199351
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1666199351
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1666199351
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1666199351
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1666199351
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1666199351
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1666199351
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1666199351
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1666199351
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1666199351
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1666199351
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1666199351
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1666199351
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1666199351
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1666199351
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1666199351
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666199351
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1666199351
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666199351
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666199351
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666199351
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666199351
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666199351
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1666199351
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666199351
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1666199351
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1666199351
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1666199351
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1666199351
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1666199351
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1666199351
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1666199351
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1666199351
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1666199351
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1666199351
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1666199351
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1666199351
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1666199351
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1666199351
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1666199351
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1666199351
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1666199351
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1666199351
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1666199351
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1666199351
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1666199351
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1666199351
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1666199351
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1666199351
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1666199351
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1666199351
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1666199351
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1666199351
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1666199351
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1666199351
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1666199351
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1666199351
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1666199351
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1666199351
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1666199351
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1666199351
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1666199351
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1666199351
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1666199351
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1666199351
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1666199351
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1666199351
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1666199351
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1666199351
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1666199351
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_513
timestamp 1666199351
transform 1 0 48300 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666199351
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666199351
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666199351
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666199351
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1666199351
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666199351
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666199351
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666199351
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1666199351
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1666199351
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666199351
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666199351
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1666199351
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1666199351
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666199351
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1666199351
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666199351
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666199351
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1666199351
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1666199351
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1666199351
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1666199351
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1666199351
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1666199351
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1666199351
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1666199351
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1666199351
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1666199351
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1666199351
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1666199351
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1666199351
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1666199351
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1666199351
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1666199351
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1666199351
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1666199351
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1666199351
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1666199351
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1666199351
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1666199351
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1666199351
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1666199351
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1666199351
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1666199351
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1666199351
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1666199351
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1666199351
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1666199351
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1666199351
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1666199351
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1666199351
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1666199351
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1666199351
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1666199351
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1666199351
transform 1 0 47564 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_513
timestamp 1666199351
transform 1 0 48300 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666199351
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1666199351
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1666199351
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666199351
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666199351
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666199351
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666199351
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666199351
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666199351
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666199351
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1666199351
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1666199351
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1666199351
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1666199351
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1666199351
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666199351
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1666199351
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1666199351
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1666199351
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1666199351
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1666199351
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1666199351
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1666199351
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1666199351
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1666199351
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1666199351
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1666199351
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1666199351
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1666199351
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1666199351
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1666199351
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1666199351
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1666199351
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1666199351
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1666199351
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1666199351
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1666199351
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1666199351
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1666199351
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1666199351
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1666199351
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1666199351
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1666199351
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1666199351
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1666199351
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1666199351
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1666199351
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1666199351
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1666199351
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1666199351
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1666199351
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1666199351
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1666199351
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1666199351
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_513
timestamp 1666199351
transform 1 0 48300 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666199351
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666199351
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1666199351
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1666199351
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1666199351
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1666199351
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666199351
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1666199351
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1666199351
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1666199351
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1666199351
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1666199351
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666199351
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666199351
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1666199351
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1666199351
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1666199351
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666199351
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1666199351
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1666199351
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1666199351
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1666199351
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1666199351
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1666199351
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1666199351
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1666199351
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1666199351
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1666199351
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1666199351
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1666199351
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1666199351
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1666199351
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1666199351
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1666199351
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1666199351
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1666199351
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1666199351
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1666199351
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1666199351
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1666199351
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1666199351
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1666199351
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1666199351
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1666199351
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1666199351
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1666199351
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1666199351
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1666199351
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1666199351
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1666199351
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1666199351
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1666199351
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1666199351
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1666199351
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_505
timestamp 1666199351
transform 1 0 47564 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_513
timestamp 1666199351
transform 1 0 48300 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1666199351
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1666199351
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1666199351
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1666199351
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1666199351
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1666199351
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1666199351
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1666199351
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1666199351
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1666199351
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1666199351
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1666199351
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1666199351
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1666199351
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1666199351
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1666199351
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1666199351
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1666199351
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1666199351
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1666199351
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1666199351
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1666199351
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1666199351
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1666199351
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1666199351
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1666199351
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1666199351
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1666199351
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1666199351
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1666199351
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1666199351
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1666199351
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1666199351
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1666199351
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1666199351
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1666199351
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1666199351
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1666199351
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1666199351
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1666199351
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1666199351
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1666199351
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1666199351
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1666199351
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1666199351
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1666199351
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1666199351
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1666199351
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1666199351
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1666199351
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1666199351
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1666199351
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1666199351
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1666199351
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_513
timestamp 1666199351
transform 1 0 48300 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1666199351
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1666199351
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1666199351
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1666199351
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1666199351
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1666199351
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1666199351
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1666199351
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1666199351
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1666199351
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1666199351
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1666199351
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1666199351
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1666199351
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1666199351
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1666199351
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1666199351
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1666199351
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1666199351
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1666199351
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1666199351
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1666199351
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1666199351
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1666199351
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1666199351
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1666199351
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1666199351
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1666199351
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1666199351
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1666199351
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1666199351
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1666199351
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1666199351
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1666199351
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1666199351
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1666199351
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1666199351
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1666199351
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1666199351
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1666199351
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1666199351
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1666199351
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1666199351
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1666199351
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1666199351
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1666199351
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1666199351
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1666199351
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1666199351
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1666199351
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1666199351
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1666199351
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1666199351
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1666199351
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1666199351
transform 1 0 47564 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_513
timestamp 1666199351
transform 1 0 48300 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1666199351
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1666199351
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1666199351
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1666199351
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1666199351
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1666199351
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1666199351
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1666199351
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1666199351
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1666199351
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1666199351
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1666199351
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1666199351
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1666199351
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1666199351
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1666199351
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1666199351
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1666199351
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1666199351
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1666199351
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1666199351
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1666199351
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1666199351
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1666199351
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1666199351
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1666199351
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1666199351
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1666199351
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1666199351
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1666199351
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1666199351
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1666199351
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1666199351
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1666199351
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1666199351
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1666199351
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1666199351
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1666199351
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1666199351
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1666199351
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1666199351
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1666199351
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1666199351
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1666199351
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1666199351
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1666199351
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1666199351
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1666199351
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1666199351
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1666199351
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1666199351
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1666199351
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1666199351
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1666199351
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_513
timestamp 1666199351
transform 1 0 48300 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1666199351
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1666199351
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1666199351
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1666199351
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1666199351
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1666199351
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1666199351
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1666199351
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1666199351
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1666199351
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1666199351
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1666199351
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1666199351
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1666199351
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1666199351
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1666199351
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1666199351
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1666199351
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1666199351
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1666199351
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1666199351
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1666199351
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1666199351
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1666199351
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1666199351
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1666199351
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1666199351
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1666199351
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1666199351
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1666199351
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1666199351
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1666199351
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1666199351
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1666199351
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1666199351
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1666199351
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1666199351
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1666199351
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1666199351
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1666199351
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1666199351
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1666199351
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1666199351
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1666199351
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1666199351
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1666199351
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1666199351
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1666199351
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1666199351
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1666199351
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1666199351
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1666199351
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1666199351
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1666199351
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1666199351
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1666199351
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1666199351
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1666199351
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1666199351
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1666199351
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1666199351
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1666199351
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1666199351
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1666199351
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1666199351
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1666199351
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1666199351
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1666199351
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1666199351
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1666199351
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1666199351
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1666199351
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1666199351
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1666199351
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1666199351
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1666199351
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1666199351
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1666199351
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1666199351
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1666199351
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1666199351
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1666199351
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1666199351
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1666199351
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1666199351
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1666199351
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1666199351
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1666199351
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1666199351
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1666199351
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1666199351
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1666199351
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1666199351
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1666199351
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1666199351
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1666199351
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1666199351
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1666199351
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1666199351
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1666199351
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1666199351
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1666199351
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1666199351
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1666199351
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1666199351
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1666199351
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1666199351
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1666199351
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1666199351
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1666199351
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1666199351
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1666199351
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1666199351
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1666199351
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1666199351
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1666199351
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1666199351
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1666199351
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1666199351
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1666199351
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1666199351
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1666199351
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1666199351
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1666199351
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1666199351
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1666199351
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1666199351
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1666199351
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1666199351
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1666199351
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1666199351
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1666199351
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1666199351
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1666199351
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1666199351
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1666199351
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1666199351
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1666199351
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1666199351
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1666199351
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1666199351
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1666199351
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1666199351
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1666199351
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1666199351
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1666199351
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1666199351
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1666199351
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1666199351
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1666199351
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1666199351
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1666199351
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1666199351
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1666199351
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1666199351
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1666199351
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1666199351
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1666199351
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1666199351
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1666199351
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1666199351
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1666199351
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1666199351
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1666199351
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1666199351
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1666199351
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1666199351
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1666199351
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1666199351
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1666199351
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1666199351
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1666199351
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1666199351
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1666199351
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1666199351
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1666199351
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1666199351
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1666199351
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1666199351
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1666199351
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1666199351
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1666199351
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1666199351
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1666199351
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1666199351
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1666199351
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1666199351
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1666199351
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1666199351
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1666199351
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1666199351
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1666199351
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1666199351
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1666199351
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1666199351
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1666199351
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1666199351
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1666199351
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1666199351
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1666199351
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1666199351
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1666199351
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1666199351
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1666199351
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1666199351
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1666199351
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1666199351
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1666199351
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1666199351
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1666199351
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1666199351
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1666199351
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1666199351
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1666199351
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1666199351
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1666199351
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1666199351
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1666199351
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1666199351
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1666199351
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1666199351
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_513
timestamp 1666199351
transform 1 0 48300 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1666199351
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1666199351
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1666199351
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1666199351
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1666199351
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1666199351
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1666199351
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1666199351
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1666199351
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1666199351
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1666199351
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1666199351
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1666199351
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1666199351
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1666199351
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1666199351
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1666199351
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1666199351
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1666199351
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1666199351
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1666199351
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1666199351
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1666199351
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1666199351
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1666199351
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1666199351
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1666199351
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1666199351
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1666199351
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1666199351
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1666199351
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1666199351
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1666199351
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1666199351
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1666199351
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1666199351
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1666199351
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1666199351
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1666199351
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1666199351
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1666199351
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1666199351
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1666199351
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1666199351
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1666199351
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1666199351
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1666199351
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1666199351
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1666199351
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1666199351
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1666199351
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1666199351
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1666199351
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1666199351
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_505
timestamp 1666199351
transform 1 0 47564 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_513
timestamp 1666199351
transform 1 0 48300 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1666199351
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1666199351
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1666199351
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1666199351
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1666199351
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1666199351
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1666199351
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1666199351
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1666199351
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1666199351
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1666199351
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1666199351
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1666199351
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1666199351
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1666199351
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1666199351
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1666199351
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1666199351
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1666199351
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1666199351
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1666199351
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1666199351
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1666199351
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1666199351
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1666199351
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1666199351
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1666199351
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1666199351
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1666199351
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1666199351
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1666199351
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1666199351
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1666199351
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1666199351
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1666199351
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1666199351
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1666199351
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1666199351
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1666199351
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1666199351
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1666199351
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1666199351
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1666199351
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1666199351
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1666199351
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1666199351
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1666199351
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1666199351
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1666199351
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1666199351
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1666199351
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1666199351
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1666199351
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1666199351
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_513
timestamp 1666199351
transform 1 0 48300 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1666199351
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1666199351
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1666199351
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1666199351
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1666199351
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1666199351
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1666199351
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1666199351
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1666199351
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1666199351
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1666199351
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1666199351
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1666199351
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1666199351
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1666199351
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1666199351
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1666199351
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1666199351
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1666199351
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1666199351
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1666199351
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1666199351
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1666199351
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1666199351
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1666199351
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1666199351
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1666199351
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1666199351
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1666199351
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1666199351
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1666199351
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1666199351
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1666199351
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1666199351
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1666199351
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1666199351
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1666199351
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1666199351
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1666199351
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1666199351
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1666199351
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1666199351
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1666199351
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1666199351
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1666199351
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1666199351
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1666199351
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1666199351
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1666199351
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1666199351
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1666199351
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1666199351
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1666199351
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1666199351
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_505
timestamp 1666199351
transform 1 0 47564 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_513
timestamp 1666199351
transform 1 0 48300 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1666199351
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1666199351
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1666199351
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1666199351
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1666199351
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1666199351
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1666199351
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1666199351
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1666199351
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1666199351
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1666199351
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1666199351
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1666199351
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1666199351
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1666199351
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1666199351
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1666199351
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1666199351
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1666199351
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1666199351
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1666199351
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1666199351
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1666199351
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1666199351
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1666199351
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1666199351
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1666199351
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1666199351
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1666199351
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1666199351
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1666199351
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1666199351
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1666199351
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1666199351
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1666199351
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1666199351
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1666199351
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1666199351
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1666199351
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1666199351
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1666199351
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1666199351
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1666199351
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1666199351
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1666199351
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1666199351
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1666199351
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1666199351
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1666199351
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1666199351
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1666199351
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1666199351
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1666199351
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1666199351
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_513
timestamp 1666199351
transform 1 0 48300 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1666199351
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1666199351
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1666199351
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1666199351
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1666199351
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1666199351
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1666199351
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1666199351
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1666199351
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1666199351
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1666199351
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1666199351
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1666199351
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1666199351
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1666199351
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1666199351
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1666199351
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1666199351
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1666199351
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1666199351
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1666199351
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1666199351
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1666199351
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1666199351
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1666199351
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1666199351
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1666199351
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1666199351
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1666199351
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1666199351
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1666199351
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1666199351
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1666199351
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1666199351
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1666199351
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1666199351
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1666199351
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1666199351
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1666199351
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1666199351
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1666199351
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1666199351
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1666199351
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1666199351
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1666199351
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1666199351
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1666199351
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1666199351
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1666199351
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1666199351
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1666199351
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1666199351
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1666199351
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1666199351
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_505
timestamp 1666199351
transform 1 0 47564 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_513
timestamp 1666199351
transform 1 0 48300 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1666199351
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1666199351
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1666199351
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1666199351
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1666199351
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1666199351
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1666199351
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1666199351
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1666199351
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1666199351
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1666199351
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1666199351
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1666199351
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1666199351
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1666199351
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1666199351
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1666199351
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1666199351
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1666199351
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1666199351
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1666199351
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1666199351
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1666199351
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1666199351
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1666199351
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1666199351
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1666199351
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1666199351
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1666199351
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1666199351
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_289
timestamp 1666199351
transform 1 0 27692 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_297
timestamp 1666199351
transform 1 0 28428 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_70_302
timestamp 1666199351
transform 1 0 28888 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1666199351
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1666199351
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1666199351
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1666199351
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1666199351
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1666199351
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1666199351
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1666199351
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1666199351
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1666199351
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1666199351
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1666199351
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1666199351
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1666199351
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1666199351
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1666199351
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1666199351
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1666199351
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1666199351
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1666199351
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1666199351
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_513
timestamp 1666199351
transform 1 0 48300 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1666199351
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1666199351
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1666199351
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1666199351
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1666199351
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1666199351
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1666199351
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1666199351
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1666199351
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1666199351
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1666199351
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1666199351
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1666199351
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1666199351
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1666199351
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1666199351
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1666199351
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1666199351
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1666199351
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1666199351
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1666199351
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1666199351
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1666199351
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1666199351
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1666199351
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1666199351
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_249
timestamp 1666199351
transform 1 0 24012 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_257
timestamp 1666199351
transform 1 0 24748 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_260
timestamp 1666199351
transform 1 0 25024 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_266
timestamp 1666199351
transform 1 0 25576 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_272
timestamp 1666199351
transform 1 0 26128 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_278
timestamp 1666199351
transform 1 0 26680 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_281
timestamp 1666199351
transform 1 0 26956 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_285
timestamp 1666199351
transform 1 0 27324 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_291
timestamp 1666199351
transform 1 0 27876 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_297
timestamp 1666199351
transform 1 0 28428 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_300
timestamp 1666199351
transform 1 0 28704 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_306
timestamp 1666199351
transform 1 0 29256 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_312
timestamp 1666199351
transform 1 0 29808 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_324
timestamp 1666199351
transform 1 0 30912 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1666199351
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1666199351
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1666199351
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1666199351
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1666199351
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1666199351
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1666199351
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1666199351
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1666199351
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1666199351
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1666199351
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1666199351
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1666199351
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1666199351
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1666199351
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1666199351
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1666199351
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1666199351
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_505
timestamp 1666199351
transform 1 0 47564 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_513
timestamp 1666199351
transform 1 0 48300 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1666199351
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1666199351
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1666199351
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1666199351
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1666199351
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1666199351
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1666199351
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1666199351
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1666199351
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1666199351
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1666199351
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1666199351
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1666199351
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1666199351
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1666199351
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1666199351
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1666199351
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1666199351
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1666199351
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1666199351
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1666199351
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1666199351
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1666199351
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1666199351
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1666199351
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1666199351
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1666199351
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_253
timestamp 1666199351
transform 1 0 24380 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_259
timestamp 1666199351
transform 1 0 24932 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_262
timestamp 1666199351
transform 1 0 25208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_266
timestamp 1666199351
transform 1 0 25576 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_289
timestamp 1666199351
transform 1 0 27692 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_295
timestamp 1666199351
transform 1 0 28244 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_299
timestamp 1666199351
transform 1 0 28612 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_303
timestamp 1666199351
transform 1 0 28980 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1666199351
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_309
timestamp 1666199351
transform 1 0 29532 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_324
timestamp 1666199351
transform 1 0 30912 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_330
timestamp 1666199351
transform 1 0 31464 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_342
timestamp 1666199351
transform 1 0 32568 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_354
timestamp 1666199351
transform 1 0 33672 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_358
timestamp 1666199351
transform 1 0 34040 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_361
timestamp 1666199351
transform 1 0 34316 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_365
timestamp 1666199351
transform 1 0 34684 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_369
timestamp 1666199351
transform 1 0 35052 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_381
timestamp 1666199351
transform 1 0 36156 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_393
timestamp 1666199351
transform 1 0 37260 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_405
timestamp 1666199351
transform 1 0 38364 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_417
timestamp 1666199351
transform 1 0 39468 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1666199351
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1666199351
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1666199351
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1666199351
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1666199351
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1666199351
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1666199351
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1666199351
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1666199351
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_513
timestamp 1666199351
transform 1 0 48300 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1666199351
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1666199351
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1666199351
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1666199351
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1666199351
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1666199351
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1666199351
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1666199351
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1666199351
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1666199351
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1666199351
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1666199351
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1666199351
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1666199351
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1666199351
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1666199351
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1666199351
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1666199351
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1666199351
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1666199351
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1666199351
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1666199351
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1666199351
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1666199351
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_225
timestamp 1666199351
transform 1 0 21804 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_233
timestamp 1666199351
transform 1 0 22540 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_236
timestamp 1666199351
transform 1 0 22816 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_257
timestamp 1666199351
transform 1 0 24748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_268
timestamp 1666199351
transform 1 0 25760 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_274
timestamp 1666199351
transform 1 0 26312 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_73_281
timestamp 1666199351
transform 1 0 26956 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_287
timestamp 1666199351
transform 1 0 27508 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_310
timestamp 1666199351
transform 1 0 29624 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_316
timestamp 1666199351
transform 1 0 30176 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_322
timestamp 1666199351
transform 1 0 30728 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_328
timestamp 1666199351
transform 1 0 31280 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_334
timestamp 1666199351
transform 1 0 31832 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_337
timestamp 1666199351
transform 1 0 32108 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_341
timestamp 1666199351
transform 1 0 32476 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_351
timestamp 1666199351
transform 1 0 33396 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_357
timestamp 1666199351
transform 1 0 33948 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_361
timestamp 1666199351
transform 1 0 34316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_364
timestamp 1666199351
transform 1 0 34592 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_370
timestamp 1666199351
transform 1 0 35144 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_376
timestamp 1666199351
transform 1 0 35696 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_382
timestamp 1666199351
transform 1 0 36248 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_388
timestamp 1666199351
transform 1 0 36800 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_393
timestamp 1666199351
transform 1 0 37260 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_397
timestamp 1666199351
transform 1 0 37628 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_403
timestamp 1666199351
transform 1 0 38180 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_415
timestamp 1666199351
transform 1 0 39284 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_427
timestamp 1666199351
transform 1 0 40388 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_439
timestamp 1666199351
transform 1 0 41492 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1666199351
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1666199351
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1666199351
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1666199351
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1666199351
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1666199351
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1666199351
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_505
timestamp 1666199351
transform 1 0 47564 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_513
timestamp 1666199351
transform 1 0 48300 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1666199351
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1666199351
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1666199351
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1666199351
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1666199351
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1666199351
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1666199351
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1666199351
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1666199351
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1666199351
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1666199351
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1666199351
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1666199351
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1666199351
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1666199351
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1666199351
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1666199351
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1666199351
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1666199351
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1666199351
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1666199351
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1666199351
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1666199351
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_221
timestamp 1666199351
transform 1 0 21436 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1666199351
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1666199351
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_253
timestamp 1666199351
transform 1 0 24380 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_266
timestamp 1666199351
transform 1 0 25576 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_272
timestamp 1666199351
transform 1 0 26128 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_287
timestamp 1666199351
transform 1 0 27508 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_291
timestamp 1666199351
transform 1 0 27876 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_305
timestamp 1666199351
transform 1 0 29164 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_309
timestamp 1666199351
transform 1 0 29532 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_323
timestamp 1666199351
transform 1 0 30820 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_329
timestamp 1666199351
transform 1 0 31372 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_335
timestamp 1666199351
transform 1 0 31924 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_341
timestamp 1666199351
transform 1 0 32476 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_347
timestamp 1666199351
transform 1 0 33028 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_350
timestamp 1666199351
transform 1 0 33304 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_354
timestamp 1666199351
transform 1 0 33672 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_362
timestamp 1666199351
transform 1 0 34408 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_365
timestamp 1666199351
transform 1 0 34684 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_370
timestamp 1666199351
transform 1 0 35144 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_377
timestamp 1666199351
transform 1 0 35788 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_385
timestamp 1666199351
transform 1 0 36524 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_391
timestamp 1666199351
transform 1 0 37076 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_397
timestamp 1666199351
transform 1 0 37628 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_403
timestamp 1666199351
transform 1 0 38180 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_409
timestamp 1666199351
transform 1 0 38732 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_415
timestamp 1666199351
transform 1 0 39284 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1666199351
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1666199351
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1666199351
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1666199351
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1666199351
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1666199351
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1666199351
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1666199351
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1666199351
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1666199351
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_513
timestamp 1666199351
transform 1 0 48300 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1666199351
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1666199351
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1666199351
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1666199351
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1666199351
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1666199351
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1666199351
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1666199351
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1666199351
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1666199351
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1666199351
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1666199351
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1666199351
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1666199351
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1666199351
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1666199351
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1666199351
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1666199351
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1666199351
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1666199351
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1666199351
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_205
timestamp 1666199351
transform 1 0 19964 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_213
timestamp 1666199351
transform 1 0 20700 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_220
timestamp 1666199351
transform 1 0 21344 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_225
timestamp 1666199351
transform 1 0 21804 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_234
timestamp 1666199351
transform 1 0 22632 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_252
timestamp 1666199351
transform 1 0 24288 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_259
timestamp 1666199351
transform 1 0 24932 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_265
timestamp 1666199351
transform 1 0 25484 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_278
timestamp 1666199351
transform 1 0 26680 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_281
timestamp 1666199351
transform 1 0 26956 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_296
timestamp 1666199351
transform 1 0 28336 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_304
timestamp 1666199351
transform 1 0 29072 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_319
timestamp 1666199351
transform 1 0 30452 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_325
timestamp 1666199351
transform 1 0 31004 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_331
timestamp 1666199351
transform 1 0 31556 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1666199351
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_337
timestamp 1666199351
transform 1 0 32108 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_343
timestamp 1666199351
transform 1 0 32660 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_356
timestamp 1666199351
transform 1 0 33856 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_363
timestamp 1666199351
transform 1 0 34500 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_367
timestamp 1666199351
transform 1 0 34868 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_390
timestamp 1666199351
transform 1 0 36984 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_393
timestamp 1666199351
transform 1 0 37260 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_397
timestamp 1666199351
transform 1 0 37628 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_403
timestamp 1666199351
transform 1 0 38180 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_426
timestamp 1666199351
transform 1 0 40296 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_438
timestamp 1666199351
transform 1 0 41400 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_446
timestamp 1666199351
transform 1 0 42136 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1666199351
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1666199351
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1666199351
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1666199351
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1666199351
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1666199351
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_505
timestamp 1666199351
transform 1 0 47564 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_513
timestamp 1666199351
transform 1 0 48300 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1666199351
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1666199351
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1666199351
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1666199351
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1666199351
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1666199351
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1666199351
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1666199351
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1666199351
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1666199351
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1666199351
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1666199351
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1666199351
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1666199351
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1666199351
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1666199351
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1666199351
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1666199351
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1666199351
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1666199351
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1666199351
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_197
timestamp 1666199351
transform 1 0 19228 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_203
timestamp 1666199351
transform 1 0 19780 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_214
timestamp 1666199351
transform 1 0 20792 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_231
timestamp 1666199351
transform 1 0 22356 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_243
timestamp 1666199351
transform 1 0 23460 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_250
timestamp 1666199351
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_253
timestamp 1666199351
transform 1 0 24380 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_277
timestamp 1666199351
transform 1 0 26588 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_298
timestamp 1666199351
transform 1 0 28520 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_76_305
timestamp 1666199351
transform 1 0 29164 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_309
timestamp 1666199351
transform 1 0 29532 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_316
timestamp 1666199351
transform 1 0 30176 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_344
timestamp 1666199351
transform 1 0 32752 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_362
timestamp 1666199351
transform 1 0 34408 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_365
timestamp 1666199351
transform 1 0 34684 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_389
timestamp 1666199351
transform 1 0 36892 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_396
timestamp 1666199351
transform 1 0 37536 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_411
timestamp 1666199351
transform 1 0 38916 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_76_417
timestamp 1666199351
transform 1 0 39468 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_421
timestamp 1666199351
transform 1 0 39836 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_425
timestamp 1666199351
transform 1 0 40204 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_431
timestamp 1666199351
transform 1 0 40756 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_437
timestamp 1666199351
transform 1 0 41308 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_443
timestamp 1666199351
transform 1 0 41860 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_455
timestamp 1666199351
transform 1 0 42964 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_467
timestamp 1666199351
transform 1 0 44068 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1666199351
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1666199351
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1666199351
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1666199351
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_513
timestamp 1666199351
transform 1 0 48300 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1666199351
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1666199351
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1666199351
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1666199351
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1666199351
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1666199351
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1666199351
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1666199351
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1666199351
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1666199351
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1666199351
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1666199351
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1666199351
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1666199351
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1666199351
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1666199351
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1666199351
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1666199351
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1666199351
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_181
timestamp 1666199351
transform 1 0 17756 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_185
timestamp 1666199351
transform 1 0 18124 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_188
timestamp 1666199351
transform 1 0 18400 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_192
timestamp 1666199351
transform 1 0 18768 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_196
timestamp 1666199351
transform 1 0 19136 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_213
timestamp 1666199351
transform 1 0 20700 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_77_221
timestamp 1666199351
transform 1 0 21436 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_225
timestamp 1666199351
transform 1 0 21804 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_241
timestamp 1666199351
transform 1 0 23276 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_245
timestamp 1666199351
transform 1 0 23644 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_258
timestamp 1666199351
transform 1 0 24840 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_269
timestamp 1666199351
transform 1 0 25852 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_278
timestamp 1666199351
transform 1 0 26680 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_281
timestamp 1666199351
transform 1 0 26956 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_285
timestamp 1666199351
transform 1 0 27324 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_295
timestamp 1666199351
transform 1 0 28244 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_315
timestamp 1666199351
transform 1 0 30084 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_334
timestamp 1666199351
transform 1 0 31832 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_337
timestamp 1666199351
transform 1 0 32108 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_347
timestamp 1666199351
transform 1 0 33028 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_353
timestamp 1666199351
transform 1 0 33580 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_364
timestamp 1666199351
transform 1 0 34592 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_370
timestamp 1666199351
transform 1 0 35144 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_387
timestamp 1666199351
transform 1 0 36708 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1666199351
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_393
timestamp 1666199351
transform 1 0 37260 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_407
timestamp 1666199351
transform 1 0 38548 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_420
timestamp 1666199351
transform 1 0 39744 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_433
timestamp 1666199351
transform 1 0 40940 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_439
timestamp 1666199351
transform 1 0 41492 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_77_445
timestamp 1666199351
transform 1 0 42044 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_449
timestamp 1666199351
transform 1 0 42412 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_453
timestamp 1666199351
transform 1 0 42780 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_465
timestamp 1666199351
transform 1 0 43884 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_477
timestamp 1666199351
transform 1 0 44988 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_489
timestamp 1666199351
transform 1 0 46092 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_501
timestamp 1666199351
transform 1 0 47196 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_505
timestamp 1666199351
transform 1 0 47564 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_513
timestamp 1666199351
transform 1 0 48300 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1666199351
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1666199351
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1666199351
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1666199351
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1666199351
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1666199351
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1666199351
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1666199351
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1666199351
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1666199351
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1666199351
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1666199351
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1666199351
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1666199351
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1666199351
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1666199351
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1666199351
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1666199351
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_177
timestamp 1666199351
transform 1 0 17388 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1666199351
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1666199351
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_197
timestamp 1666199351
transform 1 0 19228 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_201
timestamp 1666199351
transform 1 0 19596 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_215
timestamp 1666199351
transform 1 0 20884 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_230
timestamp 1666199351
transform 1 0 22264 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_243
timestamp 1666199351
transform 1 0 23460 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_250
timestamp 1666199351
transform 1 0 24104 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_78_253
timestamp 1666199351
transform 1 0 24380 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_260
timestamp 1666199351
transform 1 0 25024 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_276
timestamp 1666199351
transform 1 0 26496 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_282
timestamp 1666199351
transform 1 0 27048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_295
timestamp 1666199351
transform 1 0 28244 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_303
timestamp 1666199351
transform 1 0 28980 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1666199351
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_309
timestamp 1666199351
transform 1 0 29532 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_322
timestamp 1666199351
transform 1 0 30728 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_340
timestamp 1666199351
transform 1 0 32384 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_355
timestamp 1666199351
transform 1 0 33764 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_362
timestamp 1666199351
transform 1 0 34408 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_365
timestamp 1666199351
transform 1 0 34684 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_380
timestamp 1666199351
transform 1 0 36064 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_396
timestamp 1666199351
transform 1 0 37536 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_418
timestamp 1666199351
transform 1 0 39560 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_421
timestamp 1666199351
transform 1 0 39836 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_426
timestamp 1666199351
transform 1 0 40296 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_442
timestamp 1666199351
transform 1 0 41768 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_448
timestamp 1666199351
transform 1 0 42320 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_454
timestamp 1666199351
transform 1 0 42872 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_460
timestamp 1666199351
transform 1 0 43424 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_472
timestamp 1666199351
transform 1 0 44528 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1666199351
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1666199351
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1666199351
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_513
timestamp 1666199351
transform 1 0 48300 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1666199351
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1666199351
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1666199351
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1666199351
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1666199351
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1666199351
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1666199351
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1666199351
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1666199351
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1666199351
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1666199351
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1666199351
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1666199351
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1666199351
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1666199351
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1666199351
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1666199351
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1666199351
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_169
timestamp 1666199351
transform 1 0 16652 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_173
timestamp 1666199351
transform 1 0 17020 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_176
timestamp 1666199351
transform 1 0 17296 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_183
timestamp 1666199351
transform 1 0 17940 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_201
timestamp 1666199351
transform 1 0 19596 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_207
timestamp 1666199351
transform 1 0 20148 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_218
timestamp 1666199351
transform 1 0 21160 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_79_225
timestamp 1666199351
transform 1 0 21804 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_231
timestamp 1666199351
transform 1 0 22356 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_248
timestamp 1666199351
transform 1 0 23920 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_254
timestamp 1666199351
transform 1 0 24472 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_272
timestamp 1666199351
transform 1 0 26128 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_278
timestamp 1666199351
transform 1 0 26680 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_281
timestamp 1666199351
transform 1 0 26956 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_285
timestamp 1666199351
transform 1 0 27324 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_301
timestamp 1666199351
transform 1 0 28796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_318
timestamp 1666199351
transform 1 0 30360 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_326
timestamp 1666199351
transform 1 0 31096 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_333
timestamp 1666199351
transform 1 0 31740 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_337
timestamp 1666199351
transform 1 0 32108 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_361
timestamp 1666199351
transform 1 0 34316 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_372
timestamp 1666199351
transform 1 0 35328 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_390
timestamp 1666199351
transform 1 0 36984 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_393
timestamp 1666199351
transform 1 0 37260 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_409
timestamp 1666199351
transform 1 0 38732 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_417
timestamp 1666199351
transform 1 0 39468 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_435
timestamp 1666199351
transform 1 0 41124 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_442
timestamp 1666199351
transform 1 0 41768 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_79_449
timestamp 1666199351
transform 1 0 42412 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_454
timestamp 1666199351
transform 1 0 42872 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_460
timestamp 1666199351
transform 1 0 43424 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_466
timestamp 1666199351
transform 1 0 43976 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_478
timestamp 1666199351
transform 1 0 45080 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_490
timestamp 1666199351
transform 1 0 46184 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_502
timestamp 1666199351
transform 1 0 47288 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_505
timestamp 1666199351
transform 1 0 47564 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_513
timestamp 1666199351
transform 1 0 48300 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1666199351
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1666199351
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1666199351
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1666199351
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1666199351
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1666199351
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1666199351
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1666199351
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1666199351
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1666199351
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1666199351
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1666199351
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1666199351
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1666199351
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1666199351
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1666199351
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_153
timestamp 1666199351
transform 1 0 15180 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_161
timestamp 1666199351
transform 1 0 15916 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_166
timestamp 1666199351
transform 1 0 16376 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_186
timestamp 1666199351
transform 1 0 18216 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_194
timestamp 1666199351
transform 1 0 18952 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_197
timestamp 1666199351
transform 1 0 19228 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_201
timestamp 1666199351
transform 1 0 19596 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_212
timestamp 1666199351
transform 1 0 20608 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_218
timestamp 1666199351
transform 1 0 21160 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_235
timestamp 1666199351
transform 1 0 22724 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_248
timestamp 1666199351
transform 1 0 23920 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1666199351
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_267
timestamp 1666199351
transform 1 0 25668 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_287
timestamp 1666199351
transform 1 0 27508 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_293
timestamp 1666199351
transform 1 0 28060 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_306
timestamp 1666199351
transform 1 0 29256 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_309
timestamp 1666199351
transform 1 0 29532 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_320
timestamp 1666199351
transform 1 0 30544 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_327
timestamp 1666199351
transform 1 0 31188 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_331
timestamp 1666199351
transform 1 0 31556 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_348
timestamp 1666199351
transform 1 0 33120 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_359
timestamp 1666199351
transform 1 0 34132 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1666199351
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_365
timestamp 1666199351
transform 1 0 34684 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_370
timestamp 1666199351
transform 1 0 35144 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_377
timestamp 1666199351
transform 1 0 35788 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_381
timestamp 1666199351
transform 1 0 36156 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_396
timestamp 1666199351
transform 1 0 37536 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_402
timestamp 1666199351
transform 1 0 38088 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_416
timestamp 1666199351
transform 1 0 39376 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_421
timestamp 1666199351
transform 1 0 39836 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_427
timestamp 1666199351
transform 1 0 40388 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_444
timestamp 1666199351
transform 1 0 41952 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_451
timestamp 1666199351
transform 1 0 42596 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_458
timestamp 1666199351
transform 1 0 43240 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_465
timestamp 1666199351
transform 1 0 43884 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_471
timestamp 1666199351
transform 1 0 44436 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1666199351
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1666199351
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1666199351
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1666199351
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_513
timestamp 1666199351
transform 1 0 48300 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1666199351
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1666199351
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1666199351
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1666199351
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1666199351
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1666199351
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_57
timestamp 1666199351
transform 1 0 6348 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_64
timestamp 1666199351
transform 1 0 6992 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_76
timestamp 1666199351
transform 1 0 8096 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_88
timestamp 1666199351
transform 1 0 9200 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_100
timestamp 1666199351
transform 1 0 10304 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1666199351
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1666199351
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_137
timestamp 1666199351
transform 1 0 13708 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_81_148
timestamp 1666199351
transform 1 0 14720 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_154
timestamp 1666199351
transform 1 0 15272 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_158
timestamp 1666199351
transform 1 0 15640 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_166
timestamp 1666199351
transform 1 0 16376 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_169
timestamp 1666199351
transform 1 0 16652 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_182
timestamp 1666199351
transform 1 0 17848 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_202
timestamp 1666199351
transform 1 0 19688 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_211
timestamp 1666199351
transform 1 0 20516 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_222
timestamp 1666199351
transform 1 0 21528 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_81_225
timestamp 1666199351
transform 1 0 21804 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_232
timestamp 1666199351
transform 1 0 22448 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_254
timestamp 1666199351
transform 1 0 24472 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_260
timestamp 1666199351
transform 1 0 25024 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_278
timestamp 1666199351
transform 1 0 26680 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_281
timestamp 1666199351
transform 1 0 26956 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_286
timestamp 1666199351
transform 1 0 27416 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_312
timestamp 1666199351
transform 1 0 29808 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_316
timestamp 1666199351
transform 1 0 30176 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_333
timestamp 1666199351
transform 1 0 31740 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_81_337
timestamp 1666199351
transform 1 0 32108 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_350
timestamp 1666199351
transform 1 0 33304 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_371
timestamp 1666199351
transform 1 0 35236 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_387
timestamp 1666199351
transform 1 0 36708 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1666199351
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_393
timestamp 1666199351
transform 1 0 37260 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_407
timestamp 1666199351
transform 1 0 38548 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_426
timestamp 1666199351
transform 1 0 40296 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_433
timestamp 1666199351
transform 1 0 40940 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_440
timestamp 1666199351
transform 1 0 41584 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_446
timestamp 1666199351
transform 1 0 42136 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_449
timestamp 1666199351
transform 1 0 42412 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_454
timestamp 1666199351
transform 1 0 42872 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_461
timestamp 1666199351
transform 1 0 43516 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_468
timestamp 1666199351
transform 1 0 44160 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_475
timestamp 1666199351
transform 1 0 44804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_482
timestamp 1666199351
transform 1 0 45448 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_489
timestamp 1666199351
transform 1 0 46092 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_501
timestamp 1666199351
transform 1 0 47196 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_505
timestamp 1666199351
transform 1 0 47564 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_513
timestamp 1666199351
transform 1 0 48300 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1666199351
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1666199351
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1666199351
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_29
timestamp 1666199351
transform 1 0 3772 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_40
timestamp 1666199351
transform 1 0 4784 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_47
timestamp 1666199351
transform 1 0 5428 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_54
timestamp 1666199351
transform 1 0 6072 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_57
timestamp 1666199351
transform 1 0 6348 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_66
timestamp 1666199351
transform 1 0 7176 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_73
timestamp 1666199351
transform 1 0 7820 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_80
timestamp 1666199351
transform 1 0 8464 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_85
timestamp 1666199351
transform 1 0 8924 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_90
timestamp 1666199351
transform 1 0 9384 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_96
timestamp 1666199351
transform 1 0 9936 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_100
timestamp 1666199351
transform 1 0 10304 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_106
timestamp 1666199351
transform 1 0 10856 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_110
timestamp 1666199351
transform 1 0 11224 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_113
timestamp 1666199351
transform 1 0 11500 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_124
timestamp 1666199351
transform 1 0 12512 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_132
timestamp 1666199351
transform 1 0 13248 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_136
timestamp 1666199351
transform 1 0 13616 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_141
timestamp 1666199351
transform 1 0 14076 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_152
timestamp 1666199351
transform 1 0 15088 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_159
timestamp 1666199351
transform 1 0 15732 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_166
timestamp 1666199351
transform 1 0 16376 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_169
timestamp 1666199351
transform 1 0 16652 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_179
timestamp 1666199351
transform 1 0 17572 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_190
timestamp 1666199351
transform 1 0 18584 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_82_197
timestamp 1666199351
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_206
timestamp 1666199351
transform 1 0 20056 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_214
timestamp 1666199351
transform 1 0 20792 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_222
timestamp 1666199351
transform 1 0 21528 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_225
timestamp 1666199351
transform 1 0 21804 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_234
timestamp 1666199351
transform 1 0 22632 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_243
timestamp 1666199351
transform 1 0 23460 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1666199351
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_253
timestamp 1666199351
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_267
timestamp 1666199351
transform 1 0 25668 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_274
timestamp 1666199351
transform 1 0 26312 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_82_281
timestamp 1666199351
transform 1 0 26956 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_295
timestamp 1666199351
transform 1 0 28244 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_301
timestamp 1666199351
transform 1 0 28796 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_306
timestamp 1666199351
transform 1 0 29256 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1666199351
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_313
timestamp 1666199351
transform 1 0 29900 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_329
timestamp 1666199351
transform 1 0 31372 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_335
timestamp 1666199351
transform 1 0 31924 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_337
timestamp 1666199351
transform 1 0 32108 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_355
timestamp 1666199351
transform 1 0 33764 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_362
timestamp 1666199351
transform 1 0 34408 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_365
timestamp 1666199351
transform 1 0 34684 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_379
timestamp 1666199351
transform 1 0 35972 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_386
timestamp 1666199351
transform 1 0 36616 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_82_393
timestamp 1666199351
transform 1 0 37260 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_398
timestamp 1666199351
transform 1 0 37720 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_406
timestamp 1666199351
transform 1 0 38456 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_414
timestamp 1666199351
transform 1 0 39192 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_82_421
timestamp 1666199351
transform 1 0 39836 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_427
timestamp 1666199351
transform 1 0 40388 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_433
timestamp 1666199351
transform 1 0 40940 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_441
timestamp 1666199351
transform 1 0 41676 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_447
timestamp 1666199351
transform 1 0 42228 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_449
timestamp 1666199351
transform 1 0 42412 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_454
timestamp 1666199351
transform 1 0 42872 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_461
timestamp 1666199351
transform 1 0 43516 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_468
timestamp 1666199351
transform 1 0 44160 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_474
timestamp 1666199351
transform 1 0 44712 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1666199351
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_482
timestamp 1666199351
transform 1 0 45448 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_489
timestamp 1666199351
transform 1 0 46092 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_496
timestamp 1666199351
transform 1 0 46736 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_505
timestamp 1666199351
transform 1 0 47564 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_513
timestamp 1666199351
transform 1 0 48300 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666199351
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666199351
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666199351
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666199351
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666199351
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666199351
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666199351
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666199351
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666199351
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666199351
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666199351
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666199351
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666199351
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666199351
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666199351
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666199351
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666199351
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666199351
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666199351
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666199351
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666199351
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666199351
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666199351
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666199351
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666199351
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666199351
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666199351
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666199351
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666199351
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666199351
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666199351
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666199351
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666199351
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666199351
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666199351
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666199351
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666199351
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666199351
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666199351
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666199351
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666199351
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666199351
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666199351
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666199351
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666199351
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666199351
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666199351
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666199351
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666199351
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666199351
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666199351
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666199351
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666199351
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666199351
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666199351
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666199351
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666199351
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666199351
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666199351
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666199351
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666199351
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666199351
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666199351
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666199351
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666199351
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666199351
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666199351
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666199351
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666199351
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666199351
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666199351
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666199351
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666199351
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666199351
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666199351
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666199351
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666199351
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666199351
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666199351
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666199351
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666199351
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666199351
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666199351
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666199351
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666199351
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666199351
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666199351
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666199351
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666199351
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666199351
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666199351
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666199351
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666199351
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666199351
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666199351
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666199351
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666199351
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666199351
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666199351
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666199351
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666199351
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666199351
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666199351
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666199351
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666199351
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666199351
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666199351
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666199351
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666199351
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666199351
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666199351
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666199351
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666199351
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666199351
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666199351
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666199351
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666199351
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666199351
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666199351
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666199351
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666199351
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666199351
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666199351
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666199351
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666199351
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666199351
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666199351
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666199351
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666199351
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666199351
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666199351
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666199351
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666199351
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666199351
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666199351
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666199351
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666199351
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666199351
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1666199351
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1666199351
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1666199351
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1666199351
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1666199351
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1666199351
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1666199351
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1666199351
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1666199351
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1666199351
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1666199351
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1666199351
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1666199351
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1666199351
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1666199351
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1666199351
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1666199351
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1666199351
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1666199351
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1666199351
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1666199351
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1666199351
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1666199351
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1666199351
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1666199351
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1666199351
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1666199351
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1666199351
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666199351
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666199351
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666199351
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666199351
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666199351
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666199351
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666199351
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666199351
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666199351
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666199351
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666199351
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666199351
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666199351
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666199351
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666199351
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666199351
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666199351
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666199351
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666199351
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666199351
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666199351
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666199351
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666199351
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666199351
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666199351
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666199351
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666199351
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666199351
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666199351
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666199351
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666199351
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666199351
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666199351
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666199351
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666199351
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666199351
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666199351
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666199351
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666199351
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666199351
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666199351
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666199351
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666199351
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666199351
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666199351
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666199351
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666199351
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666199351
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666199351
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666199351
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666199351
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666199351
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666199351
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666199351
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666199351
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666199351
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666199351
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666199351
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666199351
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666199351
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666199351
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666199351
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666199351
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666199351
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666199351
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666199351
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666199351
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666199351
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666199351
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666199351
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666199351
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666199351
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666199351
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666199351
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666199351
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666199351
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666199351
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666199351
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666199351
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666199351
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666199351
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666199351
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666199351
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666199351
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666199351
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666199351
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666199351
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666199351
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666199351
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666199351
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666199351
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666199351
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666199351
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666199351
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666199351
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666199351
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666199351
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666199351
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666199351
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666199351
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666199351
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666199351
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666199351
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666199351
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666199351
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666199351
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666199351
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666199351
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666199351
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666199351
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666199351
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666199351
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666199351
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666199351
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666199351
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666199351
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666199351
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666199351
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666199351
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666199351
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666199351
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666199351
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666199351
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666199351
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666199351
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666199351
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666199351
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666199351
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666199351
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666199351
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666199351
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666199351
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666199351
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666199351
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666199351
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666199351
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666199351
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666199351
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666199351
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666199351
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666199351
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666199351
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666199351
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666199351
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666199351
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666199351
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666199351
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666199351
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666199351
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666199351
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666199351
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666199351
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666199351
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666199351
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666199351
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666199351
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666199351
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666199351
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666199351
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666199351
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666199351
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666199351
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666199351
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666199351
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666199351
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666199351
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666199351
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666199351
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666199351
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666199351
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666199351
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666199351
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666199351
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666199351
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666199351
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666199351
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666199351
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666199351
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666199351
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666199351
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666199351
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666199351
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666199351
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666199351
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666199351
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666199351
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666199351
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666199351
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666199351
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666199351
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666199351
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666199351
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666199351
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666199351
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666199351
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666199351
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666199351
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666199351
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666199351
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666199351
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666199351
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666199351
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666199351
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666199351
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666199351
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666199351
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666199351
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666199351
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666199351
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666199351
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666199351
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666199351
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666199351
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666199351
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666199351
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666199351
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666199351
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666199351
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666199351
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666199351
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666199351
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666199351
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666199351
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666199351
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666199351
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666199351
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666199351
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666199351
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666199351
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666199351
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666199351
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666199351
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666199351
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666199351
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666199351
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666199351
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666199351
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666199351
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666199351
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666199351
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666199351
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666199351
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666199351
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666199351
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666199351
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666199351
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666199351
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666199351
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666199351
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666199351
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666199351
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666199351
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666199351
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666199351
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666199351
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666199351
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666199351
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666199351
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666199351
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666199351
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666199351
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666199351
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666199351
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666199351
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666199351
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666199351
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666199351
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666199351
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666199351
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666199351
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666199351
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666199351
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666199351
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666199351
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666199351
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666199351
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666199351
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666199351
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666199351
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666199351
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666199351
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666199351
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666199351
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666199351
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666199351
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666199351
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666199351
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666199351
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666199351
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666199351
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666199351
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666199351
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666199351
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666199351
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666199351
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666199351
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666199351
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666199351
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666199351
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666199351
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666199351
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666199351
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666199351
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666199351
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666199351
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666199351
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666199351
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666199351
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666199351
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666199351
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666199351
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666199351
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666199351
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666199351
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666199351
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666199351
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666199351
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666199351
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666199351
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666199351
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666199351
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666199351
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666199351
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666199351
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666199351
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666199351
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666199351
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666199351
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666199351
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666199351
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666199351
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666199351
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666199351
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666199351
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666199351
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666199351
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666199351
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666199351
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666199351
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666199351
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666199351
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666199351
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666199351
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666199351
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666199351
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666199351
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666199351
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666199351
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666199351
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666199351
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666199351
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666199351
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666199351
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666199351
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666199351
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666199351
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666199351
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666199351
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666199351
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666199351
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666199351
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666199351
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666199351
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666199351
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666199351
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666199351
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666199351
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666199351
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666199351
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666199351
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666199351
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666199351
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666199351
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666199351
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666199351
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666199351
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666199351
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666199351
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666199351
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666199351
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666199351
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666199351
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666199351
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666199351
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666199351
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666199351
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666199351
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666199351
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666199351
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666199351
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666199351
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666199351
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666199351
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666199351
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666199351
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666199351
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666199351
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666199351
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666199351
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666199351
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666199351
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666199351
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666199351
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666199351
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666199351
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666199351
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666199351
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666199351
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666199351
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666199351
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666199351
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666199351
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666199351
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666199351
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666199351
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666199351
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666199351
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666199351
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666199351
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666199351
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666199351
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666199351
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666199351
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666199351
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666199351
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666199351
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666199351
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666199351
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666199351
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666199351
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666199351
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666199351
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666199351
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666199351
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666199351
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666199351
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666199351
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666199351
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666199351
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666199351
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666199351
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666199351
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666199351
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666199351
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666199351
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666199351
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666199351
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666199351
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666199351
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666199351
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666199351
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666199351
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666199351
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666199351
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666199351
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666199351
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666199351
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666199351
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666199351
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666199351
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666199351
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666199351
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666199351
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666199351
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666199351
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666199351
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666199351
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666199351
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666199351
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666199351
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666199351
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666199351
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666199351
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666199351
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666199351
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666199351
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666199351
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666199351
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666199351
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666199351
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666199351
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666199351
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666199351
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666199351
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666199351
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666199351
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666199351
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666199351
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666199351
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666199351
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666199351
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666199351
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666199351
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666199351
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666199351
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666199351
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666199351
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666199351
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666199351
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666199351
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666199351
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666199351
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666199351
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666199351
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666199351
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666199351
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666199351
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666199351
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666199351
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666199351
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666199351
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666199351
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666199351
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666199351
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666199351
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666199351
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666199351
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666199351
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666199351
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666199351
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666199351
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666199351
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666199351
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666199351
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666199351
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666199351
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666199351
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666199351
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666199351
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666199351
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666199351
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666199351
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666199351
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666199351
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666199351
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666199351
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666199351
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666199351
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666199351
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666199351
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666199351
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666199351
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666199351
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666199351
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666199351
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666199351
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666199351
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666199351
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666199351
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666199351
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666199351
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666199351
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666199351
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666199351
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666199351
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666199351
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666199351
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666199351
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666199351
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666199351
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666199351
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666199351
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666199351
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666199351
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666199351
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666199351
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666199351
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666199351
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666199351
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666199351
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666199351
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666199351
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666199351
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666199351
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666199351
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666199351
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666199351
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666199351
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666199351
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666199351
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666199351
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666199351
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666199351
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666199351
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666199351
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666199351
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666199351
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666199351
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666199351
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666199351
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666199351
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666199351
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666199351
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666199351
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666199351
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666199351
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666199351
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666199351
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666199351
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666199351
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666199351
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666199351
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666199351
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666199351
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666199351
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666199351
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666199351
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666199351
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666199351
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666199351
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666199351
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666199351
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666199351
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666199351
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666199351
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666199351
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666199351
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666199351
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666199351
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666199351
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666199351
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666199351
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666199351
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666199351
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666199351
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666199351
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666199351
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666199351
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666199351
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666199351
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666199351
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666199351
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666199351
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666199351
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666199351
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666199351
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666199351
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666199351
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666199351
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666199351
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666199351
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666199351
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666199351
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666199351
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666199351
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666199351
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666199351
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666199351
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666199351
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666199351
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666199351
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666199351
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666199351
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666199351
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666199351
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666199351
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666199351
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666199351
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666199351
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666199351
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666199351
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666199351
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666199351
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666199351
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666199351
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666199351
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666199351
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666199351
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666199351
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666199351
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666199351
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666199351
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666199351
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666199351
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666199351
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666199351
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666199351
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666199351
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666199351
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666199351
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666199351
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666199351
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666199351
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666199351
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666199351
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666199351
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666199351
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666199351
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666199351
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666199351
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666199351
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666199351
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666199351
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666199351
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666199351
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666199351
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666199351
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666199351
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666199351
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666199351
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666199351
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666199351
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666199351
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666199351
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666199351
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666199351
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666199351
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666199351
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666199351
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666199351
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666199351
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666199351
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666199351
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666199351
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666199351
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666199351
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666199351
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666199351
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666199351
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666199351
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666199351
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666199351
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666199351
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666199351
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666199351
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666199351
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666199351
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666199351
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666199351
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666199351
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666199351
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666199351
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666199351
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666199351
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666199351
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666199351
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666199351
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666199351
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666199351
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666199351
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666199351
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666199351
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666199351
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666199351
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666199351
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666199351
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666199351
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666199351
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666199351
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666199351
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666199351
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666199351
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666199351
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666199351
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666199351
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666199351
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666199351
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666199351
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666199351
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666199351
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666199351
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666199351
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666199351
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666199351
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _170_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 20516 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _171_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 20424 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _172_
timestamp 1666199351
transform 1 0 20700 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _173_
timestamp 1666199351
transform 1 0 26404 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_4  _174_
timestamp 1666199351
transform -1 0 30728 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _175_
timestamp 1666199351
transform -1 0 30176 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _176_
timestamp 1666199351
transform 1 0 28796 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _177_
timestamp 1666199351
transform -1 0 29164 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _178_
timestamp 1666199351
transform -1 0 30176 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _179_
timestamp 1666199351
transform 1 0 26220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_4  _180_
timestamp 1666199351
transform 1 0 27324 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _181_
timestamp 1666199351
transform -1 0 28612 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _182_
timestamp 1666199351
transform 1 0 26220 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _183_
timestamp 1666199351
transform 1 0 26404 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _184_
timestamp 1666199351
transform 1 0 26220 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _185_
timestamp 1666199351
transform -1 0 25668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_4  _186_
timestamp 1666199351
transform -1 0 26036 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _187_
timestamp 1666199351
transform 1 0 25392 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _188_
timestamp 1666199351
transform -1 0 25760 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _189_
timestamp 1666199351
transform 1 0 25116 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _190_
timestamp 1666199351
transform 1 0 23644 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _191_
timestamp 1666199351
transform -1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_4  _192_
timestamp 1666199351
transform 1 0 24564 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _193_
timestamp 1666199351
transform -1 0 25024 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _194_
timestamp 1666199351
transform 1 0 23644 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _195_
timestamp 1666199351
transform 1 0 21068 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _196_
timestamp 1666199351
transform 1 0 22816 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _197_
timestamp 1666199351
transform 1 0 21436 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_4  _198_
timestamp 1666199351
transform 1 0 22632 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _199_
timestamp 1666199351
transform -1 0 22908 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _200_
timestamp 1666199351
transform 1 0 21620 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _201_
timestamp 1666199351
transform 1 0 21068 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _202_
timestamp 1666199351
transform 1 0 21528 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _203_
timestamp 1666199351
transform 1 0 19504 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_4  _204_
timestamp 1666199351
transform 1 0 21068 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _205_
timestamp 1666199351
transform 1 0 20240 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _206_
timestamp 1666199351
transform 1 0 20240 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _207_
timestamp 1666199351
transform -1 0 20240 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _208_
timestamp 1666199351
transform -1 0 20424 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _209_
timestamp 1666199351
transform -1 0 21160 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _210_
timestamp 1666199351
transform -1 0 31096 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_4  _211_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 29716 0 1 44608
box -38 -48 1050 592
use sky130_fd_sc_hd__o31a_4  _212_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 29164 0 -1 43520
box -38 -48 1326 592
use sky130_fd_sc_hd__xnor2_4  _213_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 26588 0 1 43520
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_4  _214_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 22264 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_4  _215_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 29716 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_4  _216_
timestamp 1666199351
transform -1 0 29624 0 -1 42432
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_4  _217_
timestamp 1666199351
transform -1 0 25760 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _218_
timestamp 1666199351
transform 1 0 28888 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_4  _219_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 28612 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__a21bo_4  _220_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 29164 0 -1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_4  _221_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 27692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__or2b_4  _222_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 29716 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _223_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 29256 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _224_
timestamp 1666199351
transform 1 0 27140 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _225_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 21988 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _226_
timestamp 1666199351
transform -1 0 25576 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _227_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 23000 0 -1 43520
box -38 -48 1326 592
use sky130_fd_sc_hd__a21oi_4  _228_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 27968 0 1 42432
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _229_
timestamp 1666199351
transform -1 0 22356 0 1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _230_
timestamp 1666199351
transform 1 0 24656 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_4  _231_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 23276 0 -1 44608
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_4  _232_
timestamp 1666199351
transform -1 0 20792 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _233_
timestamp 1666199351
transform -1 0 39192 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_4  _234_
timestamp 1666199351
transform -1 0 40296 0 -1 46784
box -38 -48 1050 592
use sky130_fd_sc_hd__o31a_4  _235_
timestamp 1666199351
transform 1 0 35696 0 -1 45696
box -38 -48 1326 592
use sky130_fd_sc_hd__xnor2_4  _236_
timestamp 1666199351
transform 1 0 32292 0 -1 45696
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_4  _237_
timestamp 1666199351
transform -1 0 34132 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_4  _238_
timestamp 1666199351
transform 1 0 36432 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_4  _239_
timestamp 1666199351
transform -1 0 36984 0 -1 43520
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_4  _240_
timestamp 1666199351
transform -1 0 34592 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _241_
timestamp 1666199351
transform 1 0 39100 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_4  _242_
timestamp 1666199351
transform 1 0 38088 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__a21bo_4  _243_
timestamp 1666199351
transform 1 0 38180 0 1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_4  _244_
timestamp 1666199351
transform 1 0 37628 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__or2b_4  _245_
timestamp 1666199351
transform -1 0 40940 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _246_
timestamp 1666199351
transform -1 0 38916 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _247_
timestamp 1666199351
transform 1 0 37444 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _248_
timestamp 1666199351
transform -1 0 33764 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _249_
timestamp 1666199351
transform -1 0 34408 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _250_
timestamp 1666199351
transform 1 0 33120 0 1 43520
box -38 -48 1326 592
use sky130_fd_sc_hd__a21oi_4  _251_
timestamp 1666199351
transform 1 0 35512 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _252_
timestamp 1666199351
transform -1 0 31832 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _253_
timestamp 1666199351
transform -1 0 41676 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_4  _254_
timestamp 1666199351
transform -1 0 32384 0 1 44608
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_4  _255_
timestamp 1666199351
transform -1 0 21160 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_4  _256_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 19688 0 1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_4  _257_
timestamp 1666199351
transform 1 0 19504 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__o22a_4  _258_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 18308 0 -1 45696
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_4  _259_
timestamp 1666199351
transform -1 0 26680 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_4  _260_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 26036 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__o21a_4  _261_
timestamp 1666199351
transform 1 0 27140 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_4  _262_
timestamp 1666199351
transform -1 0 26680 0 -1 46784
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_4  _263_
timestamp 1666199351
transform -1 0 40940 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_4  _264_
timestamp 1666199351
transform 1 0 40480 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__o21a_4  _265_
timestamp 1666199351
transform 1 0 40664 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_4  _266_
timestamp 1666199351
transform -1 0 41124 0 -1 45696
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _267_
timestamp 1666199351
transform -1 0 18952 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _268_
timestamp 1666199351
transform -1 0 17848 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _269_
timestamp 1666199351
transform -1 0 16376 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _270_
timestamp 1666199351
transform 1 0 19964 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _271_
timestamp 1666199351
transform 1 0 21068 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_4  _272_
timestamp 1666199351
transform -1 0 18216 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__or2b_4  _273_
timestamp 1666199351
transform 1 0 27416 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _274_
timestamp 1666199351
transform -1 0 29808 0 -1 46784
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _275_
timestamp 1666199351
transform -1 0 28980 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _276_
timestamp 1666199351
transform 1 0 25392 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _277_
timestamp 1666199351
transform 1 0 24840 0 -1 45696
box -38 -48 1326 592
use sky130_fd_sc_hd__o21a_4  _278_
timestamp 1666199351
transform 1 0 24564 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__or2b_4  _279_
timestamp 1666199351
transform 1 0 38916 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _280_
timestamp 1666199351
transform -1 0 40296 0 -1 43520
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _281_
timestamp 1666199351
transform -1 0 38456 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _282_
timestamp 1666199351
transform 1 0 37444 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _283_
timestamp 1666199351
transform 1 0 36248 0 1 45696
box -38 -48 1326 592
use sky130_fd_sc_hd__o21a_4  _284_
timestamp 1666199351
transform 1 0 35604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _285_
timestamp 1666199351
transform -1 0 18584 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _286_
timestamp 1666199351
transform 1 0 18124 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _287_
timestamp 1666199351
transform -1 0 20056 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _288_
timestamp 1666199351
transform -1 0 17572 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_4  _289_
timestamp 1666199351
transform 1 0 18216 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__a21o_4  _290_
timestamp 1666199351
transform -1 0 26680 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _291_
timestamp 1666199351
transform 1 0 25208 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _292_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 25668 0 1 41344
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_4  _293_
timestamp 1666199351
transform 1 0 26864 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _294_
timestamp 1666199351
transform -1 0 28336 0 -1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__a32o_4  _295_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 26956 0 1 43520
box -38 -48 1602 592
use sky130_fd_sc_hd__a21o_4  _296_
timestamp 1666199351
transform 1 0 34868 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _297_
timestamp 1666199351
transform -1 0 33304 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _298_
timestamp 1666199351
transform -1 0 36892 0 1 43520
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_4  _299_
timestamp 1666199351
transform -1 0 35328 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _300_
timestamp 1666199351
transform 1 0 34868 0 1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__a32o_4  _301_
timestamp 1666199351
transform 1 0 33672 0 -1 46784
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_4  _302_
timestamp 1666199351
transform 1 0 21988 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _303_
timestamp 1666199351
transform -1 0 21528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _304_
timestamp 1666199351
transform -1 0 21528 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _305_
timestamp 1666199351
transform 1 0 22080 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_4  _306_
timestamp 1666199351
transform -1 0 22724 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__a21oi_4  _307_
timestamp 1666199351
transform 1 0 23552 0 -1 42432
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_4  _308_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 22724 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_4  _309_
timestamp 1666199351
transform 1 0 21620 0 1 42432
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_4  _310_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 23920 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _311_
timestamp 1666199351
transform 1 0 23736 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _312_
timestamp 1666199351
transform 1 0 24564 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _313_
timestamp 1666199351
transform 1 0 22632 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _314_
timestamp 1666199351
transform 1 0 32752 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_4  _315_
timestamp 1666199351
transform 1 0 32292 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_4  _316_
timestamp 1666199351
transform -1 0 32752 0 1 43520
box -38 -48 2062 592
use sky130_fd_sc_hd__o21a_4  _317_
timestamp 1666199351
transform 1 0 32660 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__a211oi_4  _318_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 33120 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__a21o_4  _319_
timestamp 1666199351
transform 1 0 30268 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__a211oi_4  _320_
timestamp 1666199351
transform -1 0 31740 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__o221a_4  _321_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 22448 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__o32a_4  _322_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 24472 0 -1 46784
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  _323_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 41584 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _324_
timestamp 1666199351
transform -1 0 42872 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _325_
timestamp 1666199351
transform -1 0 40296 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _326_
timestamp 1666199351
transform -1 0 42872 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _327_
timestamp 1666199351
transform -1 0 43516 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _328_
timestamp 1666199351
transform -1 0 43240 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _329_
timestamp 1666199351
transform -1 0 42872 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _330_
timestamp 1666199351
transform -1 0 44804 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _331_
timestamp 1666199351
transform -1 0 46092 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _332_
timestamp 1666199351
transform -1 0 46092 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _333_
timestamp 1666199351
transform 1 0 5796 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _334_
timestamp 1666199351
transform 1 0 6900 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _335_
timestamp 1666199351
transform 1 0 8188 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _336_
timestamp 1666199351
transform 1 0 23828 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _337_
timestamp 1666199351
transform -1 0 26312 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _338_
timestamp 1666199351
transform 1 0 23184 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _339_
timestamp 1666199351
transform -1 0 29164 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _340_
timestamp 1666199351
transform -1 0 34408 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _341_
timestamp 1666199351
transform -1 0 36616 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _342_
timestamp 1666199351
transform -1 0 35788 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _343_
timestamp 1666199351
transform -1 0 34408 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _344_
timestamp 1666199351
transform -1 0 40940 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _345_
timestamp 1666199351
transform -1 0 35788 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _346_
timestamp 1666199351
transform -1 0 37536 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _347_
timestamp 1666199351
transform -1 0 43516 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _348_
timestamp 1666199351
transform -1 0 41768 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _349_
timestamp 1666199351
transform -1 0 42596 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _350_
timestamp 1666199351
transform -1 0 44160 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _351_
timestamp 1666199351
transform -1 0 44160 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _352_
timestamp 1666199351
transform -1 0 43884 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _353_
timestamp 1666199351
transform -1 0 45448 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _354_
timestamp 1666199351
transform -1 0 45448 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _355_
timestamp 1666199351
transform -1 0 46736 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _356_
timestamp 1666199351
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _357_
timestamp 1666199351
transform 1 0 12144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _358_
timestamp 1666199351
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _359_
timestamp 1666199351
transform 1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _360_
timestamp 1666199351
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _361_
timestamp 1666199351
transform 1 0 13432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _362_
timestamp 1666199351
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _363_
timestamp 1666199351
transform 1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _364_
timestamp 1666199351
transform 1 0 13524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _365_
timestamp 1666199351
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _366_
timestamp 1666199351
transform 1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _367_
timestamp 1666199351
transform 1 0 14168 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _368_
timestamp 1666199351
transform 1 0 13524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _369_
timestamp 1666199351
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _370_
timestamp 1666199351
transform 1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _371_
timestamp 1666199351
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _372_
timestamp 1666199351
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _373_
timestamp 1666199351
transform 1 0 16100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _374_
timestamp 1666199351
transform 1 0 17020 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _375_
timestamp 1666199351
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _376_
timestamp 1666199351
transform 1 0 16744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _377_
timestamp 1666199351
transform 1 0 16100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _378_
timestamp 1666199351
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _379_
timestamp 1666199351
transform 1 0 17664 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _380_
timestamp 1666199351
transform 1 0 16100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _381_
timestamp 1666199351
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _382_
timestamp 1666199351
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _383_
timestamp 1666199351
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _384_
timestamp 1666199351
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _385_
timestamp 1666199351
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _386_
timestamp 1666199351
transform 1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _387_
timestamp 1666199351
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _388_
timestamp 1666199351
transform -1 0 30636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _389_
timestamp 1666199351
transform -1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _390_
timestamp 1666199351
transform -1 0 31280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _391_
timestamp 1666199351
transform -1 0 32568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _392_
timestamp 1666199351
transform -1 0 31924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _393_
timestamp 1666199351
transform -1 0 32568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _394_
timestamp 1666199351
transform -1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _395_
timestamp 1666199351
transform -1 0 32568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _396_
timestamp 1666199351
transform -1 0 33856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _397_
timestamp 1666199351
transform -1 0 33212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _398_
timestamp 1666199351
transform -1 0 33212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _399_
timestamp 1666199351
transform -1 0 33856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _400_
timestamp 1666199351
transform -1 0 33856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _401_
timestamp 1666199351
transform -1 0 35144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _402_
timestamp 1666199351
transform -1 0 34500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _403_
timestamp 1666199351
transform -1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _404_
timestamp 1666199351
transform -1 0 35144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _405_
timestamp 1666199351
transform -1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _406_
timestamp 1666199351
transform -1 0 35788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _407_
timestamp 1666199351
transform 1 0 34960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _408_
timestamp 1666199351
transform -1 0 35880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _409_
timestamp 1666199351
transform -1 0 36432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _410_
timestamp 1666199351
transform -1 0 37720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _411_
timestamp 1666199351
transform -1 0 36524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _412_
timestamp 1666199351
transform -1 0 38364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _413_
timestamp 1666199351
transform -1 0 37720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _414_
timestamp 1666199351
transform 1 0 36892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _415_
timestamp 1666199351
transform -1 0 39008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _416_
timestamp 1666199351
transform -1 0 38364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _417_
timestamp 1666199351
transform 1 0 37720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _418_
timestamp 1666199351
transform -1 0 39008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _419_
timestamp 1666199351
transform -1 0 40296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _420_
timestamp 1666199351
transform -1 0 39652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _421_
timestamp 1666199351
transform 1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _422_
timestamp 1666199351
transform -1 0 40940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _423_
timestamp 1666199351
transform -1 0 40296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _424_
timestamp 1666199351
transform -1 0 41584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _425_
timestamp 1666199351
transform -1 0 40940 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _426_
timestamp 1666199351
transform 1 0 40204 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _427_
timestamp 1666199351
transform -1 0 41584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _428_
timestamp 1666199351
transform -1 0 41124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _429_
timestamp 1666199351
transform -1 0 42872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _430_
timestamp 1666199351
transform -1 0 41768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _431_
timestamp 1666199351
transform -1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _432_
timestamp 1666199351
transform -1 0 42872 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _433_
timestamp 1666199351
transform -1 0 44160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _434_
timestamp 1666199351
transform -1 0 43516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _435_
timestamp 1666199351
transform 1 0 42688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _436_
timestamp 1666199351
transform -1 0 43608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _437_
timestamp 1666199351
transform -1 0 44160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _438_
timestamp 1666199351
transform -1 0 45448 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _439_
timestamp 1666199351
transform -1 0 44804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _440_
timestamp 1666199351
transform -1 0 46092 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _441_
timestamp 1666199351
transform -1 0 45448 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _442_
timestamp 1666199351
transform -1 0 45448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _443_
timestamp 1666199351
transform -1 0 46736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _444_
timestamp 1666199351
transform -1 0 46092 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _445_
timestamp 1666199351
transform -1 0 46092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _446_
timestamp 1666199351
transform -1 0 46736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _447_
timestamp 1666199351
transform -1 0 48024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _448_
timestamp 1666199351
transform -1 0 46736 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _449_
timestamp 1666199351
transform -1 0 47380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _450_
timestamp 1666199351
transform -1 0 48024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _451_
timestamp 1666199351
transform -1 0 48024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _455_
timestamp 1666199351
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _456_
timestamp 1666199351
transform 1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _457_
timestamp 1666199351
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _458_
timestamp 1666199351
transform 1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _459_
timestamp 1666199351
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _460_
timestamp 1666199351
transform 1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _461_
timestamp 1666199351
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _462_
timestamp 1666199351
transform 1 0 4968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _463_
timestamp 1666199351
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _464_
timestamp 1666199351
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _465_
timestamp 1666199351
transform 1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _466_
timestamp 1666199351
transform 1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _467_
timestamp 1666199351
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _468_
timestamp 1666199351
transform 1 0 6624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _469_
timestamp 1666199351
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _470_
timestamp 1666199351
transform 1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _471_
timestamp 1666199351
transform 1 0 7452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _472_
timestamp 1666199351
transform 1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _473_
timestamp 1666199351
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _474_
timestamp 1666199351
transform 1 0 8280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _475_
timestamp 1666199351
transform 1 0 7728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _476_
timestamp 1666199351
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _477_
timestamp 1666199351
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _478_
timestamp 1666199351
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _479_
timestamp 1666199351
transform 1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _480_
timestamp 1666199351
transform 1 0 9936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _481_
timestamp 1666199351
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _482_
timestamp 1666199351
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _483_
timestamp 1666199351
transform 1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _484_
timestamp 1666199351
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _485_
timestamp 1666199351
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _486_
timestamp 1666199351
transform 1 0 11500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _487_
timestamp 1666199351
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _488_
timestamp 1666199351
transform 1 0 19688 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _489_
timestamp 1666199351
transform 1 0 18676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _490_
timestamp 1666199351
transform 1 0 18032 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _491_
timestamp 1666199351
transform 1 0 19044 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _492_
timestamp 1666199351
transform 1 0 18952 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _493_
timestamp 1666199351
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _494_
timestamp 1666199351
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _495_
timestamp 1666199351
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _496_
timestamp 1666199351
transform 1 0 18676 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _497_
timestamp 1666199351
transform 1 0 21988 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _498_
timestamp 1666199351
transform 1 0 22724 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _499_
timestamp 1666199351
transform 1 0 19596 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _500_
timestamp 1666199351
transform 1 0 19320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _501_
timestamp 1666199351
transform 1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _502_
timestamp 1666199351
transform 1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _503_
timestamp 1666199351
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _504_
timestamp 1666199351
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _505_
timestamp 1666199351
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _506_
timestamp 1666199351
transform -1 0 26680 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _507_
timestamp 1666199351
transform -1 0 27416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _508_
timestamp 1666199351
transform -1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _509_
timestamp 1666199351
transform -1 0 29808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _510_
timestamp 1666199351
transform -1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _511_
timestamp 1666199351
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _512_
timestamp 1666199351
transform 1 0 27232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _513_
timestamp 1666199351
transform -1 0 28060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _514_
timestamp 1666199351
transform -1 0 29992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _515_
timestamp 1666199351
transform -1 0 30452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _516_
timestamp 1666199351
transform 1 0 28980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _517_
timestamp 1666199351
transform -1 0 30820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _518_
timestamp 1666199351
transform -1 0 31464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _519_
timestamp 1666199351
transform 1 0 28704 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _520_
timestamp 1666199351
transform 1 0 4508 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _521_
timestamp 1666199351
transform 1 0 5152 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _522_
timestamp 1666199351
transform 1 0 6716 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _523_
timestamp 1666199351
transform 1 0 7544 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _524_
timestamp 1666199351
transform -1 0 9384 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _525_
timestamp 1666199351
transform 1 0 10028 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _526_
timestamp 1666199351
transform 1 0 10948 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _527_
timestamp 1666199351
transform 1 0 12236 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _528_
timestamp 1666199351
transform 1 0 13340 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _529_
timestamp 1666199351
transform 1 0 14444 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _530_
timestamp 1666199351
transform 1 0 15364 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _531_
timestamp 1666199351
transform 1 0 14812 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _532_
timestamp 1666199351
transform 1 0 17664 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _533_
timestamp 1666199351
transform 1 0 18860 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _534_
timestamp 1666199351
transform 1 0 15456 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _535_
timestamp 1666199351
transform 1 0 21068 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _536_
timestamp 1666199351
transform 1 0 16100 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _537_
timestamp 1666199351
transform -1 0 24932 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _538_
timestamp 1666199351
transform 1 0 23828 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _539_
timestamp 1666199351
transform 1 0 23828 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _540_
timestamp 1666199351
transform -1 0 27416 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _541_
timestamp 1666199351
transform -1 0 31188 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _542_
timestamp 1666199351
transform -1 0 31740 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _543_
timestamp 1666199351
transform 1 0 29900 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _544_
timestamp 1666199351
transform -1 0 35144 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _545_
timestamp 1666199351
transform -1 0 37720 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _546_
timestamp 1666199351
transform -1 0 34500 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _547_
timestamp 1666199351
transform -1 0 35144 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _548_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 20332 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _549_
timestamp 1666199351
transform 1 0 19964 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _550_
timestamp 1666199351
transform 1 0 19688 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _551_
timestamp 1666199351
transform 1 0 21068 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _552_
timestamp 1666199351
transform 1 0 21988 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _553_
timestamp 1666199351
transform 1 0 21988 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _554_
timestamp 1666199351
transform 1 0 22356 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _555_
timestamp 1666199351
transform 1 0 22632 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _556_
timestamp 1666199351
transform 1 0 22448 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _557_
timestamp 1666199351
transform 1 0 22356 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _558_
timestamp 1666199351
transform 1 0 22908 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _559_
timestamp 1666199351
transform 1 0 23552 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _560_
timestamp 1666199351
transform 1 0 23644 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _561_
timestamp 1666199351
transform 1 0 24104 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _562_
timestamp 1666199351
transform 1 0 23920 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _563_
timestamp 1666199351
transform -1 0 25116 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _564_
timestamp 1666199351
transform 1 0 24840 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _565_
timestamp 1666199351
transform 1 0 25208 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _566_
timestamp 1666199351
transform 1 0 25208 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _567_
timestamp 1666199351
transform 1 0 25484 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _568_
timestamp 1666199351
transform 1 0 25484 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _569_
timestamp 1666199351
transform -1 0 28336 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _570_
timestamp 1666199351
transform -1 0 28336 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _571_
timestamp 1666199351
transform 1 0 27140 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _572_
timestamp 1666199351
transform -1 0 28428 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _573_
timestamp 1666199351
transform 1 0 27600 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _574_
timestamp 1666199351
transform -1 0 28796 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _575_
timestamp 1666199351
transform -1 0 28980 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _576_
timestamp 1666199351
transform -1 0 29900 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _577_
timestamp 1666199351
transform -1 0 29256 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _578_
timestamp 1666199351
transform -1 0 29900 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _579_
timestamp 1666199351
transform 1 0 29716 0 1 41344
box -38 -48 1234 592
<< labels >>
flabel metal2 s 3974 49200 4030 50000 0 FreeSans 224 90 0 0 io_active
port 0 nsew signal input
flabel metal2 s 4342 49200 4398 50000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 15382 49200 15438 50000 0 FreeSans 224 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s 16486 49200 16542 50000 0 FreeSans 224 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal2 s 17590 49200 17646 50000 0 FreeSans 224 90 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 18694 49200 18750 50000 0 FreeSans 224 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 19798 49200 19854 50000 0 FreeSans 224 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal2 s 20902 49200 20958 50000 0 FreeSans 224 90 0 0 io_in[15]
port 7 nsew signal input
flabel metal2 s 22006 49200 22062 50000 0 FreeSans 224 90 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 23110 49200 23166 50000 0 FreeSans 224 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 24214 49200 24270 50000 0 FreeSans 224 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 25318 49200 25374 50000 0 FreeSans 224 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal2 s 5446 49200 5502 50000 0 FreeSans 224 90 0 0 io_in[1]
port 12 nsew signal input
flabel metal2 s 26422 49200 26478 50000 0 FreeSans 224 90 0 0 io_in[20]
port 13 nsew signal input
flabel metal2 s 27526 49200 27582 50000 0 FreeSans 224 90 0 0 io_in[21]
port 14 nsew signal input
flabel metal2 s 28630 49200 28686 50000 0 FreeSans 224 90 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 29734 49200 29790 50000 0 FreeSans 224 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 30838 49200 30894 50000 0 FreeSans 224 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 31942 49200 31998 50000 0 FreeSans 224 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 33046 49200 33102 50000 0 FreeSans 224 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal2 s 34150 49200 34206 50000 0 FreeSans 224 90 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 35254 49200 35310 50000 0 FreeSans 224 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 36358 49200 36414 50000 0 FreeSans 224 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 6550 49200 6606 50000 0 FreeSans 224 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal2 s 37462 49200 37518 50000 0 FreeSans 224 90 0 0 io_in[30]
port 24 nsew signal input
flabel metal2 s 38566 49200 38622 50000 0 FreeSans 224 90 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 39670 49200 39726 50000 0 FreeSans 224 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal2 s 40774 49200 40830 50000 0 FreeSans 224 90 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 41878 49200 41934 50000 0 FreeSans 224 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 42982 49200 43038 50000 0 FreeSans 224 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal2 s 44086 49200 44142 50000 0 FreeSans 224 90 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 45190 49200 45246 50000 0 FreeSans 224 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 7654 49200 7710 50000 0 FreeSans 224 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal2 s 8758 49200 8814 50000 0 FreeSans 224 90 0 0 io_in[4]
port 33 nsew signal input
flabel metal2 s 9862 49200 9918 50000 0 FreeSans 224 90 0 0 io_in[5]
port 34 nsew signal input
flabel metal2 s 10966 49200 11022 50000 0 FreeSans 224 90 0 0 io_in[6]
port 35 nsew signal input
flabel metal2 s 12070 49200 12126 50000 0 FreeSans 224 90 0 0 io_in[7]
port 36 nsew signal input
flabel metal2 s 13174 49200 13230 50000 0 FreeSans 224 90 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 14278 49200 14334 50000 0 FreeSans 224 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 4710 49200 4766 50000 0 FreeSans 224 90 0 0 io_oeb[0]
port 39 nsew signal tristate
flabel metal2 s 15750 49200 15806 50000 0 FreeSans 224 90 0 0 io_oeb[10]
port 40 nsew signal tristate
flabel metal2 s 16854 49200 16910 50000 0 FreeSans 224 90 0 0 io_oeb[11]
port 41 nsew signal tristate
flabel metal2 s 17958 49200 18014 50000 0 FreeSans 224 90 0 0 io_oeb[12]
port 42 nsew signal tristate
flabel metal2 s 19062 49200 19118 50000 0 FreeSans 224 90 0 0 io_oeb[13]
port 43 nsew signal tristate
flabel metal2 s 20166 49200 20222 50000 0 FreeSans 224 90 0 0 io_oeb[14]
port 44 nsew signal tristate
flabel metal2 s 21270 49200 21326 50000 0 FreeSans 224 90 0 0 io_oeb[15]
port 45 nsew signal tristate
flabel metal2 s 22374 49200 22430 50000 0 FreeSans 224 90 0 0 io_oeb[16]
port 46 nsew signal tristate
flabel metal2 s 23478 49200 23534 50000 0 FreeSans 224 90 0 0 io_oeb[17]
port 47 nsew signal tristate
flabel metal2 s 24582 49200 24638 50000 0 FreeSans 224 90 0 0 io_oeb[18]
port 48 nsew signal tristate
flabel metal2 s 25686 49200 25742 50000 0 FreeSans 224 90 0 0 io_oeb[19]
port 49 nsew signal tristate
flabel metal2 s 5814 49200 5870 50000 0 FreeSans 224 90 0 0 io_oeb[1]
port 50 nsew signal tristate
flabel metal2 s 26790 49200 26846 50000 0 FreeSans 224 90 0 0 io_oeb[20]
port 51 nsew signal tristate
flabel metal2 s 27894 49200 27950 50000 0 FreeSans 224 90 0 0 io_oeb[21]
port 52 nsew signal tristate
flabel metal2 s 28998 49200 29054 50000 0 FreeSans 224 90 0 0 io_oeb[22]
port 53 nsew signal tristate
flabel metal2 s 30102 49200 30158 50000 0 FreeSans 224 90 0 0 io_oeb[23]
port 54 nsew signal tristate
flabel metal2 s 31206 49200 31262 50000 0 FreeSans 224 90 0 0 io_oeb[24]
port 55 nsew signal tristate
flabel metal2 s 32310 49200 32366 50000 0 FreeSans 224 90 0 0 io_oeb[25]
port 56 nsew signal tristate
flabel metal2 s 33414 49200 33470 50000 0 FreeSans 224 90 0 0 io_oeb[26]
port 57 nsew signal tristate
flabel metal2 s 34518 49200 34574 50000 0 FreeSans 224 90 0 0 io_oeb[27]
port 58 nsew signal tristate
flabel metal2 s 35622 49200 35678 50000 0 FreeSans 224 90 0 0 io_oeb[28]
port 59 nsew signal tristate
flabel metal2 s 36726 49200 36782 50000 0 FreeSans 224 90 0 0 io_oeb[29]
port 60 nsew signal tristate
flabel metal2 s 6918 49200 6974 50000 0 FreeSans 224 90 0 0 io_oeb[2]
port 61 nsew signal tristate
flabel metal2 s 37830 49200 37886 50000 0 FreeSans 224 90 0 0 io_oeb[30]
port 62 nsew signal tristate
flabel metal2 s 38934 49200 38990 50000 0 FreeSans 224 90 0 0 io_oeb[31]
port 63 nsew signal tristate
flabel metal2 s 40038 49200 40094 50000 0 FreeSans 224 90 0 0 io_oeb[32]
port 64 nsew signal tristate
flabel metal2 s 41142 49200 41198 50000 0 FreeSans 224 90 0 0 io_oeb[33]
port 65 nsew signal tristate
flabel metal2 s 42246 49200 42302 50000 0 FreeSans 224 90 0 0 io_oeb[34]
port 66 nsew signal tristate
flabel metal2 s 43350 49200 43406 50000 0 FreeSans 224 90 0 0 io_oeb[35]
port 67 nsew signal tristate
flabel metal2 s 44454 49200 44510 50000 0 FreeSans 224 90 0 0 io_oeb[36]
port 68 nsew signal tristate
flabel metal2 s 45558 49200 45614 50000 0 FreeSans 224 90 0 0 io_oeb[37]
port 69 nsew signal tristate
flabel metal2 s 8022 49200 8078 50000 0 FreeSans 224 90 0 0 io_oeb[3]
port 70 nsew signal tristate
flabel metal2 s 9126 49200 9182 50000 0 FreeSans 224 90 0 0 io_oeb[4]
port 71 nsew signal tristate
flabel metal2 s 10230 49200 10286 50000 0 FreeSans 224 90 0 0 io_oeb[5]
port 72 nsew signal tristate
flabel metal2 s 11334 49200 11390 50000 0 FreeSans 224 90 0 0 io_oeb[6]
port 73 nsew signal tristate
flabel metal2 s 12438 49200 12494 50000 0 FreeSans 224 90 0 0 io_oeb[7]
port 74 nsew signal tristate
flabel metal2 s 13542 49200 13598 50000 0 FreeSans 224 90 0 0 io_oeb[8]
port 75 nsew signal tristate
flabel metal2 s 14646 49200 14702 50000 0 FreeSans 224 90 0 0 io_oeb[9]
port 76 nsew signal tristate
flabel metal2 s 5078 49200 5134 50000 0 FreeSans 224 90 0 0 io_out[0]
port 77 nsew signal tristate
flabel metal2 s 16118 49200 16174 50000 0 FreeSans 224 90 0 0 io_out[10]
port 78 nsew signal tristate
flabel metal2 s 17222 49200 17278 50000 0 FreeSans 224 90 0 0 io_out[11]
port 79 nsew signal tristate
flabel metal2 s 18326 49200 18382 50000 0 FreeSans 224 90 0 0 io_out[12]
port 80 nsew signal tristate
flabel metal2 s 19430 49200 19486 50000 0 FreeSans 224 90 0 0 io_out[13]
port 81 nsew signal tristate
flabel metal2 s 20534 49200 20590 50000 0 FreeSans 224 90 0 0 io_out[14]
port 82 nsew signal tristate
flabel metal2 s 21638 49200 21694 50000 0 FreeSans 224 90 0 0 io_out[15]
port 83 nsew signal tristate
flabel metal2 s 22742 49200 22798 50000 0 FreeSans 224 90 0 0 io_out[16]
port 84 nsew signal tristate
flabel metal2 s 23846 49200 23902 50000 0 FreeSans 224 90 0 0 io_out[17]
port 85 nsew signal tristate
flabel metal2 s 24950 49200 25006 50000 0 FreeSans 224 90 0 0 io_out[18]
port 86 nsew signal tristate
flabel metal2 s 26054 49200 26110 50000 0 FreeSans 224 90 0 0 io_out[19]
port 87 nsew signal tristate
flabel metal2 s 6182 49200 6238 50000 0 FreeSans 224 90 0 0 io_out[1]
port 88 nsew signal tristate
flabel metal2 s 27158 49200 27214 50000 0 FreeSans 224 90 0 0 io_out[20]
port 89 nsew signal tristate
flabel metal2 s 28262 49200 28318 50000 0 FreeSans 224 90 0 0 io_out[21]
port 90 nsew signal tristate
flabel metal2 s 29366 49200 29422 50000 0 FreeSans 224 90 0 0 io_out[22]
port 91 nsew signal tristate
flabel metal2 s 30470 49200 30526 50000 0 FreeSans 224 90 0 0 io_out[23]
port 92 nsew signal tristate
flabel metal2 s 31574 49200 31630 50000 0 FreeSans 224 90 0 0 io_out[24]
port 93 nsew signal tristate
flabel metal2 s 32678 49200 32734 50000 0 FreeSans 224 90 0 0 io_out[25]
port 94 nsew signal tristate
flabel metal2 s 33782 49200 33838 50000 0 FreeSans 224 90 0 0 io_out[26]
port 95 nsew signal tristate
flabel metal2 s 34886 49200 34942 50000 0 FreeSans 224 90 0 0 io_out[27]
port 96 nsew signal tristate
flabel metal2 s 35990 49200 36046 50000 0 FreeSans 224 90 0 0 io_out[28]
port 97 nsew signal tristate
flabel metal2 s 37094 49200 37150 50000 0 FreeSans 224 90 0 0 io_out[29]
port 98 nsew signal tristate
flabel metal2 s 7286 49200 7342 50000 0 FreeSans 224 90 0 0 io_out[2]
port 99 nsew signal tristate
flabel metal2 s 38198 49200 38254 50000 0 FreeSans 224 90 0 0 io_out[30]
port 100 nsew signal tristate
flabel metal2 s 39302 49200 39358 50000 0 FreeSans 224 90 0 0 io_out[31]
port 101 nsew signal tristate
flabel metal2 s 40406 49200 40462 50000 0 FreeSans 224 90 0 0 io_out[32]
port 102 nsew signal tristate
flabel metal2 s 41510 49200 41566 50000 0 FreeSans 224 90 0 0 io_out[33]
port 103 nsew signal tristate
flabel metal2 s 42614 49200 42670 50000 0 FreeSans 224 90 0 0 io_out[34]
port 104 nsew signal tristate
flabel metal2 s 43718 49200 43774 50000 0 FreeSans 224 90 0 0 io_out[35]
port 105 nsew signal tristate
flabel metal2 s 44822 49200 44878 50000 0 FreeSans 224 90 0 0 io_out[36]
port 106 nsew signal tristate
flabel metal2 s 45926 49200 45982 50000 0 FreeSans 224 90 0 0 io_out[37]
port 107 nsew signal tristate
flabel metal2 s 8390 49200 8446 50000 0 FreeSans 224 90 0 0 io_out[3]
port 108 nsew signal tristate
flabel metal2 s 9494 49200 9550 50000 0 FreeSans 224 90 0 0 io_out[4]
port 109 nsew signal tristate
flabel metal2 s 10598 49200 10654 50000 0 FreeSans 224 90 0 0 io_out[5]
port 110 nsew signal tristate
flabel metal2 s 11702 49200 11758 50000 0 FreeSans 224 90 0 0 io_out[6]
port 111 nsew signal tristate
flabel metal2 s 12806 49200 12862 50000 0 FreeSans 224 90 0 0 io_out[7]
port 112 nsew signal tristate
flabel metal2 s 13910 49200 13966 50000 0 FreeSans 224 90 0 0 io_out[8]
port 113 nsew signal tristate
flabel metal2 s 15014 49200 15070 50000 0 FreeSans 224 90 0 0 io_out[9]
port 114 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 115 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 116 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 117 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 118 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 119 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 120 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 121 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 122 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 123 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 124 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 125 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 126 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 127 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 128 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 129 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 130 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 131 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 132 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 133 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 134 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 135 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 136 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 137 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 138 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 139 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 140 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 141 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 142 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 143 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 144 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 145 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 146 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 147 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 148 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 149 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 150 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 151 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 152 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 153 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 154 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 155 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 156 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 157 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 158 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 159 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 160 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 161 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 162 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 163 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 164 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 165 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 166 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 167 nsew signal input
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 168 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 169 nsew signal input
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 170 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 171 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 172 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 173 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 174 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 175 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 176 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 177 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 178 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 179 nsew signal input
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 180 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 181 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 182 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 183 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 184 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 185 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 186 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 187 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 188 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 189 nsew signal input
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 190 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 191 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 192 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 193 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 194 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 195 nsew signal input
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 196 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 197 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 198 nsew signal input
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 199 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 200 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 201 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 202 nsew signal input
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 203 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 204 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 205 nsew signal input
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 206 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 207 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 208 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 209 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 210 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 211 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 212 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 213 nsew signal input
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 214 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 215 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 216 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 217 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 218 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 219 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 220 nsew signal input
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 221 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 222 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 223 nsew signal input
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 224 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 225 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 226 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 227 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 228 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 229 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 230 nsew signal input
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 231 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 232 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 233 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 234 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 235 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 236 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 237 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 238 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 239 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 240 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 241 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 242 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 243 nsew signal tristate
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 244 nsew signal tristate
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 245 nsew signal tristate
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 246 nsew signal tristate
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 247 nsew signal tristate
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 248 nsew signal tristate
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 249 nsew signal tristate
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 250 nsew signal tristate
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 251 nsew signal tristate
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 252 nsew signal tristate
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 253 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 254 nsew signal tristate
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 255 nsew signal tristate
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 256 nsew signal tristate
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 257 nsew signal tristate
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 258 nsew signal tristate
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 259 nsew signal tristate
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 260 nsew signal tristate
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 261 nsew signal tristate
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 262 nsew signal tristate
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 263 nsew signal tristate
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 264 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 265 nsew signal tristate
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 266 nsew signal tristate
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 267 nsew signal tristate
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 268 nsew signal tristate
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 269 nsew signal tristate
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 270 nsew signal tristate
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 271 nsew signal tristate
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 272 nsew signal tristate
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 273 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 274 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 275 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 276 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 277 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 278 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 279 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 280 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 281 nsew signal tristate
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 282 nsew signal tristate
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 283 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 284 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 285 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 286 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 287 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 288 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 289 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 290 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 291 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 292 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 293 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 294 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 295 nsew signal tristate
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 296 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 297 nsew signal tristate
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 298 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 299 nsew signal tristate
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 300 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 301 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 302 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 303 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 304 nsew signal tristate
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 305 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 306 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 307 nsew signal tristate
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 308 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 309 nsew signal tristate
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 310 nsew signal tristate
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 311 nsew signal tristate
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 312 nsew signal tristate
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 313 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 314 nsew signal tristate
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 315 nsew signal tristate
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 316 nsew signal tristate
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 317 nsew signal tristate
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 318 nsew signal tristate
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 319 nsew signal tristate
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 320 nsew signal tristate
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 321 nsew signal tristate
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 322 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 323 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 324 nsew signal tristate
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 325 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 326 nsew signal tristate
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 327 nsew signal tristate
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 328 nsew signal tristate
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 329 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 330 nsew signal tristate
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 331 nsew signal tristate
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 332 nsew signal tristate
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 333 nsew signal tristate
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 334 nsew signal tristate
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 335 nsew signal tristate
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 336 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 337 nsew signal tristate
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 338 nsew signal tristate
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 339 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 340 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 341 nsew signal tristate
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 342 nsew signal tristate
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 343 nsew signal tristate
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 344 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 345 nsew signal tristate
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 346 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 347 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 348 nsew signal tristate
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 349 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 350 nsew signal tristate
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 351 nsew signal tristate
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 352 nsew signal tristate
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 353 nsew signal tristate
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 354 nsew signal tristate
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 355 nsew signal tristate
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 356 nsew signal tristate
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 357 nsew signal tristate
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 358 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 359 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 360 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 361 nsew signal tristate
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 362 nsew signal tristate
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 363 nsew signal tristate
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 364 nsew signal tristate
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 365 nsew signal tristate
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 366 nsew signal tristate
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 367 nsew signal tristate
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 368 nsew signal tristate
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 369 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 370 nsew signal tristate
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 371 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 372 nsew signal input
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 373 nsew signal input
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 374 nsew signal input
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 375 nsew signal input
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 376 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 377 nsew signal input
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 378 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 379 nsew signal input
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 380 nsew signal input
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 381 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 382 nsew signal input
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 383 nsew signal input
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 384 nsew signal input
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 385 nsew signal input
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 386 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 387 nsew signal input
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 388 nsew signal input
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 389 nsew signal input
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 390 nsew signal input
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 391 nsew signal input
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 392 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 393 nsew signal input
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 394 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 395 nsew signal input
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 396 nsew signal input
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 397 nsew signal input
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 398 nsew signal input
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 399 nsew signal input
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 400 nsew signal input
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 401 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 402 nsew signal input
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 403 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 404 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 405 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 406 nsew signal input
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 407 nsew signal input
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 408 nsew signal input
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 409 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 410 nsew signal input
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 411 nsew signal input
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 412 nsew signal input
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 413 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 414 nsew signal input
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 415 nsew signal input
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 416 nsew signal input
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 417 nsew signal input
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 418 nsew signal input
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 419 nsew signal input
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 420 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 421 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 422 nsew signal input
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 423 nsew signal input
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 424 nsew signal input
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 425 nsew signal input
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 426 nsew signal input
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 427 nsew signal input
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 428 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 429 nsew signal input
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 430 nsew signal input
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 431 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 432 nsew signal input
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 433 nsew signal input
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 434 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 435 nsew signal input
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 436 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 437 nsew signal input
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 438 nsew signal input
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 439 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 440 nsew signal input
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 441 nsew signal input
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 442 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 443 nsew signal input
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 444 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 445 nsew signal input
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 446 nsew signal input
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 447 nsew signal input
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 448 nsew signal input
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 449 nsew signal input
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 450 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 451 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 452 nsew signal input
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 453 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 454 nsew signal input
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 455 nsew signal input
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 456 nsew signal input
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 457 nsew signal input
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 458 nsew signal input
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 459 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 460 nsew signal input
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 461 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 462 nsew signal input
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 463 nsew signal input
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 464 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 465 nsew signal input
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 466 nsew signal input
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 467 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 468 nsew signal input
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 469 nsew signal input
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 470 nsew signal input
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 471 nsew signal input
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 472 nsew signal input
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 473 nsew signal input
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 474 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 475 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 476 nsew signal input
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 477 nsew signal input
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 478 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 479 nsew signal input
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 480 nsew signal input
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 481 nsew signal input
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 482 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 483 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 484 nsew signal input
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 485 nsew signal input
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 486 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 487 nsew signal input
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 488 nsew signal input
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 489 nsew signal input
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 490 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 491 nsew signal input
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 492 nsew signal input
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 493 nsew signal input
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 494 nsew signal input
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 495 nsew signal input
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 496 nsew signal input
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 497 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 498 nsew signal input
flabel metal4 s 4208 2128 4528 47376 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 34928 2128 35248 47376 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 19568 2128 19888 47376 0 FreeSans 1920 90 0 0 vssd1
port 500 nsew ground bidirectional
flabel metal2 s 2410 0 2466 800 0 FreeSans 224 90 0 0 wb_clk_i
port 501 nsew signal input
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 wb_rst_i
port 502 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 503 nsew signal tristate
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 504 nsew signal input
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 505 nsew signal input
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 506 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 507 nsew signal input
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 508 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 509 nsew signal input
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 510 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 511 nsew signal input
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 512 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 513 nsew signal input
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 514 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 515 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 516 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 517 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 518 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 519 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 520 nsew signal input
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 521 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 522 nsew signal input
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 523 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 524 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 525 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 526 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 527 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 528 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 529 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 530 nsew signal input
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 531 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 532 nsew signal input
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 533 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 534 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 535 nsew signal input
flabel metal2 s 2686 0 2742 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 536 nsew signal input
flabel metal2 s 3054 0 3110 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 537 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 538 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 539 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 540 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 541 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 542 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 543 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 544 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 545 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 546 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 547 nsew signal input
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 548 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 549 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 550 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 551 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 552 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 553 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 554 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 555 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 556 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 557 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 558 nsew signal input
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 559 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 560 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 561 nsew signal input
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 562 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 563 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 564 nsew signal input
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 565 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 566 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 567 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 568 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 569 nsew signal tristate
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 570 nsew signal tristate
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 571 nsew signal tristate
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 572 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 573 nsew signal tristate
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 574 nsew signal tristate
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 575 nsew signal tristate
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 576 nsew signal tristate
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 577 nsew signal tristate
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 578 nsew signal tristate
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 579 nsew signal tristate
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 580 nsew signal tristate
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 581 nsew signal tristate
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 582 nsew signal tristate
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 583 nsew signal tristate
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 584 nsew signal tristate
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 585 nsew signal tristate
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 586 nsew signal tristate
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 587 nsew signal tristate
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 588 nsew signal tristate
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 589 nsew signal tristate
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 590 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 591 nsew signal tristate
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 592 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 593 nsew signal tristate
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 594 nsew signal tristate
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 595 nsew signal tristate
flabel metal2 s 4894 0 4950 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 596 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 597 nsew signal tristate
flabel metal2 s 5446 0 5502 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 598 nsew signal tristate
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 599 nsew signal tristate
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 600 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 601 nsew signal input
flabel metal2 s 3606 0 3662 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 602 nsew signal input
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 603 nsew signal input
flabel metal2 s 4342 0 4398 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 604 nsew signal input
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 605 nsew signal input
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 wbs_we_i
port 606 nsew signal input
rlabel metal1 24978 47328 24978 47328 0 vccd1
rlabel metal1 24978 46784 24978 46784 0 vssd1
rlabel metal2 20378 2686 20378 2686 0 _000_
rlabel metal2 26450 45118 26450 45118 0 _001_
rlabel metal2 29762 42976 29762 42976 0 _002_
rlabel metal2 28014 43180 28014 43180 0 _003_
rlabel metal1 22770 43282 22770 43282 0 _004_
rlabel metal2 21942 44574 21942 44574 0 _005_
rlabel metal2 29486 42398 29486 42398 0 _006_
rlabel metal2 26634 41786 26634 41786 0 _007_
rlabel metal1 24748 42194 24748 42194 0 _008_
rlabel metal1 29808 45934 29808 45934 0 _009_
rlabel metal1 28566 45424 28566 45424 0 _010_
rlabel metal2 28934 45696 28934 45696 0 _011_
rlabel metal2 28014 44642 28014 44642 0 _012_
rlabel metal2 29670 46342 29670 46342 0 _013_
rlabel metal2 27646 45356 27646 45356 0 _014_
rlabel metal1 27232 43282 27232 43282 0 _015_
rlabel metal1 23092 43214 23092 43214 0 _016_
rlabel metal2 23782 42398 23782 42398 0 _017_
rlabel metal1 21482 43724 21482 43724 0 _018_
rlabel metal2 22954 43452 22954 43452 0 _019_
rlabel metal2 20562 44064 20562 44064 0 _020_
rlabel metal2 23138 44948 23138 44948 0 _021_
rlabel metal1 20378 44336 20378 44336 0 _022_
rlabel metal2 20194 44608 20194 44608 0 _023_
rlabel metal1 37352 44846 37352 44846 0 _024_
rlabel metal1 38962 44880 38962 44880 0 _025_
rlabel metal1 35328 45526 35328 45526 0 _026_
rlabel metal1 33626 44880 33626 44880 0 _027_
rlabel metal1 32200 44370 32200 44370 0 _028_
rlabel metal2 36478 44030 36478 44030 0 _029_
rlabel metal1 35926 43690 35926 43690 0 _030_
rlabel metal2 34178 43962 34178 43962 0 _031_
rlabel metal2 39330 45050 39330 45050 0 _032_
rlabel metal2 38686 44302 38686 44302 0 _033_
rlabel metal2 38594 44574 38594 44574 0 _034_
rlabel metal2 38318 44846 38318 44846 0 _035_
rlabel metal2 39974 43792 39974 43792 0 _036_
rlabel metal1 38456 43962 38456 43962 0 _037_
rlabel metal1 36892 44370 36892 44370 0 _038_
rlabel metal1 33304 44302 33304 44302 0 _039_
rlabel metal2 33810 43248 33810 43248 0 _040_
rlabel metal2 32338 44404 32338 44404 0 _041_
rlabel metal1 32430 44200 32430 44200 0 _042_
rlabel metal2 20930 45186 20930 45186 0 _043_
rlabel metal1 38686 45526 38686 45526 0 _044_
rlabel metal1 21068 45458 21068 45458 0 _045_
rlabel metal1 19964 45458 19964 45458 0 _046_
rlabel metal2 26358 45220 26358 45220 0 _047_
rlabel metal1 27508 46138 27508 46138 0 _048_
rlabel metal1 26542 46614 26542 46614 0 _049_
rlabel metal1 20158 45934 20158 45934 0 _050_
rlabel metal2 40618 46444 40618 46444 0 _051_
rlabel metal1 41354 44914 41354 44914 0 _052_
rlabel metal1 40526 44914 40526 44914 0 _053_
rlabel metal2 39882 44914 39882 44914 0 _054_
rlabel metal2 18722 46580 18722 46580 0 _055_
rlabel metal1 16790 46546 16790 46546 0 _056_
rlabel metal2 21114 45118 21114 45118 0 _057_
rlabel metal1 28658 44438 28658 44438 0 _058_
rlabel metal1 25438 47056 25438 47056 0 _059_
rlabel metal2 26082 45220 26082 45220 0 _060_
rlabel metal2 25438 45186 25438 45186 0 _061_
rlabel metal1 25024 45526 25024 45526 0 _062_
rlabel metal2 19918 47090 19918 47090 0 _063_
rlabel metal2 39422 43724 39422 43724 0 _064_
rlabel metal1 37904 43350 37904 43350 0 _065_
rlabel metal1 38226 47124 38226 47124 0 _066_
rlabel metal2 36938 46206 36938 46206 0 _067_
rlabel metal2 36386 46308 36386 46308 0 _068_
rlabel via2 35558 46563 35558 46563 0 _069_
rlabel metal2 18170 45900 18170 45900 0 _070_
rlabel metal1 17526 47056 17526 47056 0 _071_
rlabel metal1 27140 43350 27140 43350 0 _072_
rlabel metal1 27416 43758 27416 43758 0 _073_
rlabel metal1 27370 42670 27370 42670 0 _074_
rlabel metal1 27784 42738 27784 42738 0 _075_
rlabel metal2 28198 43588 28198 43588 0 _076_
rlabel metal2 21758 44948 21758 44948 0 _077_
rlabel metal2 34454 46750 34454 46750 0 _078_
rlabel metal1 33856 46546 33856 46546 0 _079_
rlabel metal2 35558 44268 35558 44268 0 _080_
rlabel metal1 34776 45526 34776 45526 0 _081_
rlabel metal1 35282 44982 35282 44982 0 _082_
rlabel metal1 33672 46614 33672 46614 0 _083_
rlabel metal1 21758 47056 21758 47056 0 _084_
rlabel metal2 22126 46427 22126 46427 0 _085_
rlabel metal2 22678 42500 22678 42500 0 _086_
rlabel metal2 23046 43146 23046 43146 0 _087_
rlabel metal2 23230 44166 23230 44166 0 _088_
rlabel metal2 24334 46274 24334 46274 0 _089_
rlabel metal1 23000 44846 23000 44846 0 _090_
rlabel metal1 22862 45492 22862 45492 0 _091_
rlabel metal1 23782 44914 23782 44914 0 _092_
rlabel metal2 32798 43554 32798 43554 0 _093_
rlabel metal2 31878 44030 31878 44030 0 _094_
rlabel metal2 31142 45220 31142 45220 0 _095_
rlabel metal2 32062 46444 32062 46444 0 _096_
rlabel metal2 30958 46274 30958 46274 0 _097_
rlabel metal1 24058 46580 24058 46580 0 _098_
rlabel metal1 19458 4590 19458 4590 0 _099_
rlabel metal2 20930 6154 20930 6154 0 _100_
rlabel metal2 29026 6154 29026 6154 0 _101_
rlabel metal1 27968 6290 27968 6290 0 _102_
rlabel metal1 25576 6766 25576 6766 0 _103_
rlabel metal2 22862 4420 22862 4420 0 _104_
rlabel metal2 21574 3264 21574 3264 0 _105_
rlabel metal2 20562 6120 20562 6120 0 _106_
rlabel metal2 20194 3298 20194 3298 0 _107_
rlabel metal1 20010 5270 20010 5270 0 _108_
rlabel metal1 21298 4488 21298 4488 0 _109_
rlabel metal1 22080 4182 22080 4182 0 _110_
rlabel metal1 21804 2618 21804 2618 0 _111_
rlabel metal1 22586 3400 22586 3400 0 _112_
rlabel metal2 22862 2584 22862 2584 0 _113_
rlabel metal2 22678 5440 22678 5440 0 _114_
rlabel metal2 22586 6120 22586 6120 0 _115_
rlabel metal1 23046 7174 23046 7174 0 _116_
rlabel metal1 23644 4182 23644 4182 0 _117_
rlabel metal1 23828 3094 23828 3094 0 _118_
rlabel metal2 24334 5440 24334 5440 0 _119_
rlabel metal2 24150 6120 24150 6120 0 _120_
rlabel metal2 24886 7208 24886 7208 0 _121_
rlabel metal2 25070 3434 25070 3434 0 _122_
rlabel metal2 25438 3230 25438 3230 0 _123_
rlabel metal2 25438 4386 25438 4386 0 _124_
rlabel metal2 25714 6120 25714 6120 0 _125_
rlabel metal2 25714 7208 25714 7208 0 _126_
rlabel metal1 27738 4182 27738 4182 0 _127_
rlabel metal2 28106 3230 28106 3230 0 _128_
rlabel metal1 27002 5270 27002 5270 0 _129_
rlabel metal2 28198 5848 28198 5848 0 _130_
rlabel metal2 27830 6562 27830 6562 0 _131_
rlabel metal1 28566 2312 28566 2312 0 _132_
rlabel metal2 28750 3672 28750 3672 0 _133_
rlabel metal2 29670 5440 29670 5440 0 _134_
rlabel metal1 29026 4488 29026 4488 0 _135_
rlabel metal1 29992 3094 29992 3094 0 _136_
rlabel metal2 20010 45594 20010 45594 0 _137_
rlabel metal1 20194 6222 20194 6222 0 _138_
rlabel metal2 18906 3230 18906 3230 0 _139_
rlabel metal2 18262 4964 18262 4964 0 _140_
rlabel metal2 21206 4828 21206 4828 0 _141_
rlabel metal1 20654 4046 20654 4046 0 _142_
rlabel metal1 19136 2618 19136 2618 0 _143_
rlabel metal1 20700 3570 20700 3570 0 _144_
rlabel metal1 21390 2482 21390 2482 0 _145_
rlabel metal1 20746 4794 20746 4794 0 _146_
rlabel metal1 22356 7174 22356 7174 0 _147_
rlabel metal1 23000 7854 23000 7854 0 _148_
rlabel metal1 21758 3978 21758 3978 0 _149_
rlabel metal1 21666 2890 21666 2890 0 _150_
rlabel metal1 22862 5066 22862 5066 0 _151_
rlabel metal2 24058 7106 24058 7106 0 _152_
rlabel metal2 24978 7650 24978 7650 0 _153_
rlabel metal1 24978 2516 24978 2516 0 _154_
rlabel metal1 22402 2414 22402 2414 0 _155_
rlabel metal1 25346 4488 25346 4488 0 _156_
rlabel metal1 25944 6222 25944 6222 0 _157_
rlabel metal1 25852 7310 25852 7310 0 _158_
rlabel metal1 28888 4046 28888 4046 0 _159_
rlabel metal1 29900 2618 29900 2618 0 _160_
rlabel metal2 27278 4964 27278 4964 0 _161_
rlabel metal1 27876 4794 27876 4794 0 _162_
rlabel metal1 27784 7174 27784 7174 0 _163_
rlabel metal1 29210 2482 29210 2482 0 _164_
rlabel metal1 29532 3570 29532 3570 0 _165_
rlabel metal2 29762 5678 29762 5678 0 _166_
rlabel metal1 29854 4658 29854 4658 0 _167_
rlabel metal2 31234 2788 31234 2788 0 _168_
rlabel metal1 29394 41650 29394 41650 0 _169_
rlabel metal1 20056 46546 20056 46546 0 active
rlabel metal2 26266 41174 26266 41174 0 io_in[18]
rlabel metal1 28980 41174 28980 41174 0 io_in[19]
rlabel metal1 27324 41242 27324 41242 0 io_in[20]
rlabel metal1 23828 41242 23828 41242 0 io_in[21]
rlabel metal2 29670 40800 29670 40800 0 io_in[22]
rlabel metal1 32062 42330 32062 42330 0 io_in[23]
rlabel metal1 30406 43282 30406 43282 0 io_in[24]
rlabel metal2 32115 49300 32115 49300 0 io_in[25]
rlabel metal1 41446 44846 41446 44846 0 io_in[26]
rlabel metal1 38502 43826 38502 43826 0 io_in[27]
rlabel metal1 36570 42330 36570 42330 0 io_in[28]
rlabel metal2 36846 46886 36846 46886 0 io_in[29]
rlabel metal1 37260 42738 37260 42738 0 io_in[30]
rlabel metal2 41170 43180 41170 43180 0 io_in[31]
rlabel metal1 36386 43316 36386 43316 0 io_in[32]
rlabel metal2 36202 44540 36202 44540 0 io_in[33]
rlabel metal1 38870 44200 38870 44200 0 io_in[34]
rlabel metal2 43010 47661 43010 47661 0 io_in[35]
rlabel metal1 42458 44506 42458 44506 0 io_in[36]
rlabel metal2 43286 44336 43286 44336 0 io_in[37]
rlabel metal2 4738 48256 4738 48256 0 io_oeb[0]
rlabel metal2 15594 47923 15594 47923 0 io_oeb[10]
rlabel metal1 15962 47226 15962 47226 0 io_oeb[11]
rlabel metal1 17940 45458 17940 45458 0 io_oeb[12]
rlabel metal2 19090 46828 19090 46828 0 io_oeb[13]
rlabel metal1 16468 47090 16468 47090 0 io_oeb[14]
rlabel metal2 21298 46284 21298 46284 0 io_oeb[15]
rlabel metal1 17434 47090 17434 47090 0 io_oeb[16]
rlabel metal1 24196 43146 24196 43146 0 io_oeb[17]
rlabel metal1 24242 43962 24242 43962 0 io_oeb[18]
rlabel metal1 24886 47226 24886 47226 0 io_oeb[19]
rlabel metal1 5612 47226 5612 47226 0 io_oeb[1]
rlabel metal1 27002 46478 27002 46478 0 io_oeb[20]
rlabel metal1 30958 45968 30958 45968 0 io_oeb[21]
rlabel metal1 31510 45526 31510 45526 0 io_oeb[22]
rlabel metal2 30130 46624 30130 46624 0 io_oeb[23]
rlabel metal1 34546 45934 34546 45934 0 io_oeb[24]
rlabel metal2 37490 46852 37490 46852 0 io_oeb[25]
rlabel metal2 33994 47396 33994 47396 0 io_oeb[26]
rlabel metal1 34822 42738 34822 42738 0 io_oeb[27]
rlabel metal1 38594 46376 38594 46376 0 io_oeb[28]
rlabel metal1 42550 47022 42550 47022 0 io_oeb[29]
rlabel metal2 6946 47916 6946 47916 0 io_oeb[2]
rlabel metal1 40020 45050 40020 45050 0 io_oeb[30]
rlabel metal1 42044 46410 42044 46410 0 io_oeb[31]
rlabel metal1 41814 46546 41814 46546 0 io_oeb[32]
rlabel metal1 42090 46070 42090 46070 0 io_oeb[33]
rlabel metal2 42642 45499 42642 45499 0 io_oeb[34]
rlabel metal1 43976 46546 43976 46546 0 io_oeb[35]
rlabel metal2 44758 48093 44758 48093 0 io_oeb[36]
rlabel metal2 45862 47923 45862 47923 0 io_oeb[37]
rlabel metal2 7774 48263 7774 48263 0 io_oeb[3]
rlabel metal2 9154 48256 9154 48256 0 io_oeb[4]
rlabel metal2 10258 48256 10258 48256 0 io_oeb[5]
rlabel metal2 11178 48263 11178 48263 0 io_oeb[6]
rlabel metal2 12466 48256 12466 48256 0 io_oeb[7]
rlabel metal2 13570 48256 13570 48256 0 io_oeb[8]
rlabel metal2 14674 47916 14674 47916 0 io_oeb[9]
rlabel metal2 4646 45465 4646 45465 0 io_out[0]
rlabel metal2 16146 47984 16146 47984 0 io_out[10]
rlabel metal1 18262 46580 18262 46580 0 io_out[11]
rlabel metal2 18630 48093 18630 48093 0 io_out[12]
rlabel metal1 19458 46444 19458 46444 0 io_out[13]
rlabel metal1 20930 44506 20930 44506 0 io_out[14]
rlabel metal1 18630 46546 18630 46546 0 io_out[15]
rlabel metal1 22540 46410 22540 46410 0 io_out[16]
rlabel metal1 23547 46546 23547 46546 0 io_out[17]
rlabel metal1 24518 45050 24518 45050 0 io_out[18]
rlabel metal2 26082 48256 26082 48256 0 io_out[19]
rlabel metal2 6026 48263 6026 48263 0 io_out[1]
rlabel metal1 23414 46988 23414 46988 0 io_out[20]
rlabel metal1 28612 43962 28612 43962 0 io_out[21]
rlabel metal1 34178 46954 34178 46954 0 io_out[22]
rlabel metal2 36386 46937 36386 46937 0 io_out[23]
rlabel metal1 34546 46002 34546 46002 0 io_out[24]
rlabel metal1 33442 46682 33442 46682 0 io_out[25]
rlabel via2 40710 46461 40710 46461 0 io_out[26]
rlabel metal1 35512 42738 35512 42738 0 io_out[27]
rlabel metal3 37214 45628 37214 45628 0 io_out[28]
rlabel metal2 43286 46869 43286 46869 0 io_out[29]
rlabel metal2 7130 48263 7130 48263 0 io_out[2]
rlabel metal2 41492 46308 41492 46308 0 io_out[30]
rlabel metal1 40848 46138 40848 46138 0 io_out[31]
rlabel metal1 42182 47226 42182 47226 0 io_out[32]
rlabel metal1 42734 46478 42734 46478 0 io_out[33]
rlabel metal1 43148 46138 43148 46138 0 io_out[34]
rlabel metal1 44712 47226 44712 47226 0 io_out[35]
rlabel metal1 45034 46546 45034 46546 0 io_out[36]
rlabel metal1 46230 47226 46230 47226 0 io_out[37]
rlabel metal2 8418 48256 8418 48256 0 io_out[3]
rlabel metal2 9522 47950 9522 47950 0 io_out[4]
rlabel metal2 10626 48086 10626 48086 0 io_out[5]
rlabel metal2 11730 47712 11730 47712 0 io_out[6]
rlabel metal2 19458 46070 19458 46070 0 io_out[7]
rlabel metal1 21068 46002 21068 46002 0 io_out[8]
rlabel metal2 15042 47848 15042 47848 0 io_out[9]
rlabel metal2 12282 1588 12282 1588 0 la_data_out[0]
rlabel metal2 39882 1588 39882 1588 0 la_data_out[100]
rlabel metal2 40158 1792 40158 1792 0 la_data_out[101]
rlabel metal2 40434 2132 40434 2132 0 la_data_out[102]
rlabel metal2 40710 1860 40710 1860 0 la_data_out[103]
rlabel metal2 40986 2132 40986 2132 0 la_data_out[104]
rlabel metal2 41262 1622 41262 1622 0 la_data_out[105]
rlabel metal2 41538 2132 41538 2132 0 la_data_out[106]
rlabel metal2 41814 1588 41814 1588 0 la_data_out[107]
rlabel metal2 42090 1792 42090 1792 0 la_data_out[108]
rlabel metal2 42366 1656 42366 1656 0 la_data_out[109]
rlabel metal2 15042 2132 15042 2132 0 la_data_out[10]
rlabel metal2 42642 1860 42642 1860 0 la_data_out[110]
rlabel metal2 42918 2132 42918 2132 0 la_data_out[111]
rlabel metal2 43194 2132 43194 2132 0 la_data_out[112]
rlabel metal2 43470 1792 43470 1792 0 la_data_out[113]
rlabel metal2 43746 1622 43746 1622 0 la_data_out[114]
rlabel metal2 44022 1792 44022 1792 0 la_data_out[115]
rlabel metal2 44298 1554 44298 1554 0 la_data_out[116]
rlabel metal2 44574 1860 44574 1860 0 la_data_out[117]
rlabel metal2 44850 2132 44850 2132 0 la_data_out[118]
rlabel metal2 45126 1656 45126 1656 0 la_data_out[119]
rlabel metal2 15318 1860 15318 1860 0 la_data_out[11]
rlabel metal2 45402 1792 45402 1792 0 la_data_out[120]
rlabel metal2 45678 2132 45678 2132 0 la_data_out[121]
rlabel metal2 45954 1792 45954 1792 0 la_data_out[122]
rlabel metal2 46230 1588 46230 1588 0 la_data_out[123]
rlabel metal2 46506 2132 46506 2132 0 la_data_out[124]
rlabel metal2 46782 2132 46782 2132 0 la_data_out[125]
rlabel metal2 47058 1792 47058 1792 0 la_data_out[126]
rlabel metal2 47334 2132 47334 2132 0 la_data_out[127]
rlabel metal2 15594 1588 15594 1588 0 la_data_out[12]
rlabel metal2 15870 1792 15870 1792 0 la_data_out[13]
rlabel metal2 16146 2336 16146 2336 0 la_data_out[14]
rlabel metal2 16422 2132 16422 2132 0 la_data_out[15]
rlabel metal2 16698 1622 16698 1622 0 la_data_out[16]
rlabel metal2 16974 1299 16974 1299 0 la_data_out[17]
rlabel metal2 17250 2336 17250 2336 0 la_data_out[18]
rlabel metal2 17526 1860 17526 1860 0 la_data_out[19]
rlabel metal2 12558 2132 12558 2132 0 la_data_out[1]
rlabel metal2 17802 2166 17802 2166 0 la_data_out[20]
rlabel metal2 18078 1826 18078 1826 0 la_data_out[21]
rlabel metal2 18354 1554 18354 1554 0 la_data_out[22]
rlabel metal2 18630 2370 18630 2370 0 la_data_out[23]
rlabel metal2 18906 1622 18906 1622 0 la_data_out[24]
rlabel metal2 19182 2200 19182 2200 0 la_data_out[25]
rlabel metal2 19458 2336 19458 2336 0 la_data_out[26]
rlabel metal2 19734 1095 19734 1095 0 la_data_out[27]
rlabel metal2 20010 1027 20010 1027 0 la_data_out[28]
rlabel metal2 20286 1656 20286 1656 0 la_data_out[29]
rlabel metal2 12834 1622 12834 1622 0 la_data_out[2]
rlabel metal2 20562 1928 20562 1928 0 la_data_out[30]
rlabel metal2 20838 1588 20838 1588 0 la_data_out[31]
rlabel metal2 21114 3492 21114 3492 0 la_data_out[32]
rlabel metal2 21390 2098 21390 2098 0 la_data_out[33]
rlabel metal2 21666 2948 21666 2948 0 la_data_out[34]
rlabel metal2 21942 1503 21942 1503 0 la_data_out[35]
rlabel metal2 22218 1435 22218 1435 0 la_data_out[36]
rlabel metal2 22494 1860 22494 1860 0 la_data_out[37]
rlabel metal2 22770 2166 22770 2166 0 la_data_out[38]
rlabel metal2 23046 1622 23046 1622 0 la_data_out[39]
rlabel metal2 13110 2132 13110 2132 0 la_data_out[3]
rlabel metal2 23322 1503 23322 1503 0 la_data_out[40]
rlabel metal2 23598 3492 23598 3492 0 la_data_out[41]
rlabel metal2 23874 3798 23874 3798 0 la_data_out[42]
rlabel metal2 24150 2404 24150 2404 0 la_data_out[43]
rlabel metal2 24426 1860 24426 1860 0 la_data_out[44]
rlabel metal2 24702 1775 24702 1775 0 la_data_out[45]
rlabel metal2 24978 3492 24978 3492 0 la_data_out[46]
rlabel metal1 24978 7310 24978 7310 0 la_data_out[47]
rlabel metal2 25530 1622 25530 1622 0 la_data_out[48]
rlabel metal2 25806 1860 25806 1860 0 la_data_out[49]
rlabel metal2 13386 1826 13386 1826 0 la_data_out[4]
rlabel metal2 26082 1571 26082 1571 0 la_data_out[50]
rlabel metal2 26358 3458 26358 3458 0 la_data_out[51]
rlabel metal2 26634 4036 26634 4036 0 la_data_out[52]
rlabel metal2 26910 2404 26910 2404 0 la_data_out[53]
rlabel metal2 27186 1860 27186 1860 0 la_data_out[54]
rlabel metal2 27462 1775 27462 1775 0 la_data_out[55]
rlabel metal2 27738 3254 27738 3254 0 la_data_out[56]
rlabel metal2 28014 3798 28014 3798 0 la_data_out[57]
rlabel metal2 28290 1622 28290 1622 0 la_data_out[58]
rlabel metal2 28566 2166 28566 2166 0 la_data_out[59]
rlabel metal2 13662 2132 13662 2132 0 la_data_out[5]
rlabel metal2 28842 2948 28842 2948 0 la_data_out[60]
rlabel metal2 29118 2710 29118 2710 0 la_data_out[61]
rlabel metal2 29394 1860 29394 1860 0 la_data_out[62]
rlabel metal2 29670 2098 29670 2098 0 la_data_out[63]
rlabel metal2 29946 2132 29946 2132 0 la_data_out[64]
rlabel metal2 30222 1792 30222 1792 0 la_data_out[65]
rlabel metal2 30498 2132 30498 2132 0 la_data_out[66]
rlabel metal2 30774 1588 30774 1588 0 la_data_out[67]
rlabel metal2 31050 2200 31050 2200 0 la_data_out[68]
rlabel metal2 31326 1792 31326 1792 0 la_data_out[69]
rlabel metal2 13938 1792 13938 1792 0 la_data_out[6]
rlabel metal2 31602 1622 31602 1622 0 la_data_out[70]
rlabel metal2 31878 2132 31878 2132 0 la_data_out[71]
rlabel metal2 32154 1656 32154 1656 0 la_data_out[72]
rlabel metal2 32430 1792 32430 1792 0 la_data_out[73]
rlabel metal2 32706 2132 32706 2132 0 la_data_out[74]
rlabel metal2 32982 1860 32982 1860 0 la_data_out[75]
rlabel metal2 33258 2132 33258 2132 0 la_data_out[76]
rlabel metal2 33534 1622 33534 1622 0 la_data_out[77]
rlabel metal2 33810 1792 33810 1792 0 la_data_out[78]
rlabel metal2 34086 1588 34086 1588 0 la_data_out[79]
rlabel metal2 14214 1656 14214 1656 0 la_data_out[7]
rlabel metal2 34362 1792 34362 1792 0 la_data_out[80]
rlabel metal2 34638 1656 34638 1656 0 la_data_out[81]
rlabel metal2 34914 1095 34914 1095 0 la_data_out[82]
rlabel metal2 35190 1299 35190 1299 0 la_data_out[83]
rlabel metal2 35466 2132 35466 2132 0 la_data_out[84]
rlabel metal2 35742 1792 35742 1792 0 la_data_out[85]
rlabel metal2 36018 1588 36018 1588 0 la_data_out[86]
rlabel metal2 36294 2132 36294 2132 0 la_data_out[87]
rlabel metal2 36570 1622 36570 1622 0 la_data_out[88]
rlabel metal2 36846 1792 36846 1792 0 la_data_out[89]
rlabel metal2 14490 1826 14490 1826 0 la_data_out[8]
rlabel metal2 37122 2132 37122 2132 0 la_data_out[90]
rlabel metal2 37398 1554 37398 1554 0 la_data_out[91]
rlabel metal2 37674 1792 37674 1792 0 la_data_out[92]
rlabel metal2 37950 2132 37950 2132 0 la_data_out[93]
rlabel metal2 38226 1792 38226 1792 0 la_data_out[94]
rlabel metal2 38502 1656 38502 1656 0 la_data_out[95]
rlabel metal2 38778 1860 38778 1860 0 la_data_out[96]
rlabel metal2 39054 2132 39054 2132 0 la_data_out[97]
rlabel metal2 39330 1622 39330 1622 0 la_data_out[98]
rlabel metal2 39606 1792 39606 1792 0 la_data_out[99]
rlabel metal2 14766 1622 14766 1622 0 la_data_out[9]
rlabel metal2 2622 1588 2622 1588 0 wbs_ack_o
rlabel metal2 3174 1792 3174 1792 0 wbs_dat_o[0]
rlabel metal2 6302 1826 6302 1826 0 wbs_dat_o[10]
rlabel metal2 6578 1792 6578 1792 0 wbs_dat_o[11]
rlabel metal2 6854 2132 6854 2132 0 wbs_dat_o[12]
rlabel metal2 7130 1656 7130 1656 0 wbs_dat_o[13]
rlabel metal1 6463 2414 6463 2414 0 wbs_dat_o[14]
rlabel metal2 7682 2132 7682 2132 0 wbs_dat_o[15]
rlabel metal2 7958 1860 7958 1860 0 wbs_dat_o[16]
rlabel metal2 8234 1622 8234 1622 0 wbs_dat_o[17]
rlabel metal2 8510 2132 8510 2132 0 wbs_dat_o[18]
rlabel metal2 8786 1826 8786 1826 0 wbs_dat_o[19]
rlabel metal2 3542 1622 3542 1622 0 wbs_dat_o[1]
rlabel metal2 9062 1792 9062 1792 0 wbs_dat_o[20]
rlabel metal2 9338 2132 9338 2132 0 wbs_dat_o[21]
rlabel metal2 9614 1656 9614 1656 0 wbs_dat_o[22]
rlabel metal2 9890 1860 9890 1860 0 wbs_dat_o[23]
rlabel metal2 10166 2132 10166 2132 0 wbs_dat_o[24]
rlabel metal2 10442 1622 10442 1622 0 wbs_dat_o[25]
rlabel metal2 10718 1792 10718 1792 0 wbs_dat_o[26]
rlabel metal2 10994 2132 10994 2132 0 wbs_dat_o[27]
rlabel metal2 11270 1826 11270 1826 0 wbs_dat_o[28]
rlabel metal2 11546 1656 11546 1656 0 wbs_dat_o[29]
rlabel metal2 3910 1792 3910 1792 0 wbs_dat_o[2]
rlabel metal2 11822 2132 11822 2132 0 wbs_dat_o[30]
rlabel metal2 12098 1792 12098 1792 0 wbs_dat_o[31]
rlabel metal2 4278 1656 4278 1656 0 wbs_dat_o[3]
rlabel metal2 4646 1588 4646 1588 0 wbs_dat_o[4]
rlabel metal2 4922 1826 4922 1826 0 wbs_dat_o[5]
rlabel metal2 5198 2132 5198 2132 0 wbs_dat_o[6]
rlabel metal2 5474 1860 5474 1860 0 wbs_dat_o[7]
rlabel metal2 5750 1588 5750 1588 0 wbs_dat_o[8]
rlabel metal2 6026 2132 6026 2132 0 wbs_dat_o[9]
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
