magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 98 157 366 203
rect 1 21 919 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 174 47 204 177
rect 258 47 288 177
rect 446 47 476 131
rect 518 47 548 131
rect 609 47 639 131
rect 693 47 723 131
rect 811 47 841 131
<< scpmoshvt >>
rect 79 413 109 497
rect 174 297 204 497
rect 258 297 288 497
rect 429 413 459 497
rect 523 413 553 497
rect 609 413 639 497
rect 693 413 723 497
rect 811 413 841 497
<< ndiff >>
rect 124 131 174 177
rect 27 101 79 131
rect 27 67 35 101
rect 69 67 79 101
rect 27 47 79 67
rect 109 93 174 131
rect 109 59 119 93
rect 153 59 174 93
rect 109 47 174 59
rect 204 101 258 177
rect 204 67 214 101
rect 248 67 258 101
rect 204 47 258 67
rect 288 93 340 177
rect 288 59 298 93
rect 332 59 340 93
rect 288 47 340 59
rect 394 101 446 131
rect 394 67 402 101
rect 436 67 446 101
rect 394 47 446 67
rect 476 47 518 131
rect 548 47 609 131
rect 639 47 693 131
rect 723 101 811 131
rect 723 67 767 101
rect 801 67 811 101
rect 723 47 811 67
rect 841 101 893 131
rect 841 67 851 101
rect 885 67 893 101
rect 841 47 893 67
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 413 79 443
rect 109 485 174 497
rect 109 451 119 485
rect 153 451 174 485
rect 109 413 174 451
rect 124 297 174 413
rect 204 343 258 497
rect 204 309 214 343
rect 248 309 258 343
rect 204 297 258 309
rect 288 485 429 497
rect 288 451 314 485
rect 348 451 382 485
rect 416 451 429 485
rect 288 413 429 451
rect 459 477 523 497
rect 459 443 479 477
rect 513 443 523 477
rect 459 413 523 443
rect 553 485 609 497
rect 553 451 563 485
rect 597 451 609 485
rect 553 413 609 451
rect 639 477 693 497
rect 639 443 649 477
rect 683 443 693 477
rect 639 413 693 443
rect 723 485 811 497
rect 723 451 767 485
rect 801 451 811 485
rect 723 413 811 451
rect 841 477 893 497
rect 841 443 851 477
rect 885 443 893 477
rect 841 413 893 443
rect 288 297 414 413
<< ndiffc >>
rect 35 67 69 101
rect 119 59 153 93
rect 214 67 248 101
rect 298 59 332 93
rect 402 67 436 101
rect 767 67 801 101
rect 851 67 885 101
<< pdiffc >>
rect 35 443 69 477
rect 119 451 153 485
rect 214 309 248 343
rect 314 451 348 485
rect 382 451 416 485
rect 479 443 513 477
rect 563 451 597 485
rect 649 443 683 477
rect 767 451 801 485
rect 851 443 885 477
<< poly >>
rect 79 497 109 523
rect 174 497 204 523
rect 258 497 288 523
rect 429 497 459 523
rect 523 497 553 523
rect 609 497 639 523
rect 693 497 723 523
rect 811 497 841 523
rect 79 265 109 413
rect 21 249 109 265
rect 21 215 32 249
rect 66 215 109 249
rect 21 199 109 215
rect 79 131 109 199
rect 174 265 204 297
rect 258 265 288 297
rect 429 265 459 413
rect 523 346 553 413
rect 505 330 559 346
rect 505 296 515 330
rect 549 296 559 330
rect 505 280 559 296
rect 174 249 327 265
rect 174 215 283 249
rect 317 215 327 249
rect 174 199 327 215
rect 369 249 459 265
rect 369 215 379 249
rect 413 215 459 249
rect 369 199 459 215
rect 174 177 204 199
rect 258 177 288 199
rect 385 190 459 199
rect 385 146 476 190
rect 446 131 476 146
rect 518 131 548 280
rect 609 221 639 413
rect 693 281 723 413
rect 687 265 741 281
rect 687 231 697 265
rect 731 231 741 265
rect 591 205 645 221
rect 687 215 741 231
rect 811 219 841 413
rect 591 171 601 205
rect 635 171 645 205
rect 591 155 645 171
rect 609 131 639 155
rect 693 131 723 215
rect 791 203 845 219
rect 791 169 801 203
rect 835 169 845 203
rect 791 153 845 169
rect 811 131 841 153
rect 79 21 109 47
rect 174 21 204 47
rect 258 21 288 47
rect 446 21 476 47
rect 518 21 548 47
rect 609 21 639 47
rect 693 21 723 47
rect 811 21 841 47
<< polycont >>
rect 32 215 66 249
rect 515 296 549 330
rect 283 215 317 249
rect 379 215 413 249
rect 697 231 731 265
rect 601 171 635 205
rect 801 169 835 203
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 35 477 69 493
rect 103 485 169 527
rect 103 451 119 485
rect 153 451 169 485
rect 298 485 432 527
rect 298 451 314 485
rect 348 451 382 485
rect 416 451 432 485
rect 479 477 513 493
rect 35 411 69 443
rect 547 485 615 527
rect 547 451 563 485
rect 597 451 615 485
rect 649 477 683 493
rect 479 417 513 443
rect 751 485 817 527
rect 751 451 767 485
rect 801 451 817 485
rect 851 477 903 493
rect 649 417 683 443
rect 885 443 903 477
rect 851 417 903 443
rect 35 377 385 411
rect 30 249 66 327
rect 30 215 32 249
rect 30 199 66 215
rect 100 161 134 377
rect 198 309 214 343
rect 248 309 264 343
rect 35 127 134 161
rect 35 101 69 127
rect 203 101 248 309
rect 351 265 385 377
rect 447 383 683 417
rect 717 383 903 417
rect 283 249 317 265
rect 283 161 317 215
rect 351 249 413 265
rect 351 215 379 249
rect 351 199 413 215
rect 447 161 481 383
rect 717 349 751 383
rect 515 330 751 349
rect 549 315 751 330
rect 515 280 549 296
rect 670 265 731 281
rect 283 127 481 161
rect 582 205 635 255
rect 582 171 601 205
rect 35 51 69 67
rect 103 59 119 93
rect 153 59 169 93
rect 103 17 169 59
rect 203 67 214 101
rect 402 101 436 127
rect 203 51 248 67
rect 282 59 298 93
rect 332 59 348 93
rect 282 17 348 59
rect 582 84 635 171
rect 670 231 697 265
rect 670 85 731 231
rect 765 203 835 261
rect 765 169 801 203
rect 765 153 835 169
rect 869 117 903 383
rect 767 101 817 117
rect 402 51 436 67
rect 801 67 817 101
rect 767 17 817 67
rect 851 101 903 117
rect 885 67 903 101
rect 851 51 903 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 582 85 616 119 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 765 153 799 187 0 FreeSans 200 0 0 0 B_N
port 2 nsew signal input
flabel locali s 582 153 616 187 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 214 289 248 323 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 214 153 248 187 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 674 85 708 119 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
rlabel comment s 0 0 0 0 4 and4bb_2
rlabel metal1 s 0 -48 920 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 3097452
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3089516
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 23.000 0.000 
<< end >>
