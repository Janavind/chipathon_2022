magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< pwell >>
rect 547 2026 568 2075
rect 1841 2026 1862 2075
rect 1179 1269 1189 1279
rect 547 874 568 923
rect 1841 874 1862 923
<< obsli1 >>
rect 0 0 2654 2370
<< obsm1 >>
rect 0 2304 2654 2370
rect 0 1218 66 2304
rect 94 1793 122 2276
rect 150 1821 178 2304
rect 206 1793 234 2276
rect 262 1821 290 2304
rect 318 1793 346 2276
rect 374 1821 402 2304
rect 430 1793 458 2276
rect 486 1821 514 2304
rect 542 1793 570 2276
rect 598 1821 626 2304
rect 654 1793 706 2276
rect 734 1821 762 2304
rect 790 1793 818 2276
rect 846 1821 874 2304
rect 902 1793 930 2276
rect 958 1821 986 2304
rect 1014 1793 1042 2276
rect 1070 1821 1098 2304
rect 1126 1793 1154 2276
rect 1182 1821 1210 2304
rect 1238 1793 1266 2276
rect 94 1729 1266 1793
rect 94 1246 122 1729
rect 150 1218 178 1701
rect 206 1246 234 1729
rect 262 1218 290 1701
rect 318 1246 346 1729
rect 374 1218 402 1701
rect 430 1246 458 1729
rect 486 1218 514 1701
rect 542 1246 570 1729
rect 598 1218 626 1701
rect 654 1246 706 1729
rect 734 1218 762 1701
rect 790 1246 818 1729
rect 846 1218 874 1701
rect 902 1246 930 1729
rect 958 1218 986 1701
rect 1014 1246 1042 1729
rect 1070 1218 1098 1701
rect 1126 1246 1154 1729
rect 1182 1218 1210 1701
rect 1238 1246 1266 1729
rect 1294 1218 1360 2304
rect 1388 1793 1416 2276
rect 1444 1821 1472 2304
rect 1500 1793 1528 2276
rect 1556 1821 1584 2304
rect 1612 1793 1640 2276
rect 1668 1821 1696 2304
rect 1724 1793 1752 2276
rect 1780 1821 1808 2304
rect 1836 1793 1864 2276
rect 1892 1821 1920 2304
rect 1948 1793 2000 2276
rect 2028 1821 2056 2304
rect 2084 1793 2112 2276
rect 2140 1821 2168 2304
rect 2196 1793 2224 2276
rect 2252 1821 2280 2304
rect 2308 1793 2336 2276
rect 2364 1821 2392 2304
rect 2420 1793 2448 2276
rect 2476 1821 2504 2304
rect 2532 1793 2560 2276
rect 1388 1729 2560 1793
rect 1388 1246 1416 1729
rect 1444 1218 1472 1701
rect 1500 1246 1528 1729
rect 1556 1218 1584 1701
rect 1612 1246 1640 1729
rect 1668 1218 1696 1701
rect 1724 1246 1752 1729
rect 1780 1218 1808 1701
rect 1836 1246 1864 1729
rect 1892 1218 1920 1701
rect 1948 1246 2000 1729
rect 2028 1218 2056 1701
rect 2084 1246 2112 1729
rect 2140 1218 2168 1701
rect 2196 1246 2224 1729
rect 2252 1218 2280 1701
rect 2308 1246 2336 1729
rect 2364 1218 2392 1701
rect 2420 1246 2448 1729
rect 2476 1218 2504 1701
rect 2532 1246 2560 1729
rect 2588 1218 2654 2304
rect 0 1152 2654 1218
rect 0 66 66 1152
rect 94 641 122 1124
rect 150 669 178 1152
rect 206 641 234 1124
rect 262 669 290 1152
rect 318 641 346 1124
rect 374 669 402 1152
rect 430 641 458 1124
rect 486 669 514 1152
rect 542 641 570 1124
rect 598 669 626 1152
rect 654 641 706 1124
rect 734 669 762 1152
rect 790 641 818 1124
rect 846 669 874 1152
rect 902 641 930 1124
rect 958 669 986 1152
rect 1014 641 1042 1124
rect 1070 669 1098 1152
rect 1126 641 1154 1124
rect 1182 669 1210 1152
rect 1238 641 1266 1124
rect 94 577 1266 641
rect 94 94 122 577
rect 150 66 178 549
rect 206 94 234 577
rect 262 66 290 549
rect 318 94 346 577
rect 374 66 402 549
rect 430 94 458 577
rect 486 66 514 549
rect 542 94 570 577
rect 598 66 626 549
rect 654 94 706 577
rect 734 66 762 549
rect 790 94 818 577
rect 846 66 874 549
rect 902 94 930 577
rect 958 66 986 549
rect 1014 94 1042 577
rect 1070 66 1098 549
rect 1126 94 1154 577
rect 1182 66 1210 549
rect 1238 94 1266 577
rect 1294 66 1360 1152
rect 1388 641 1416 1124
rect 1444 669 1472 1152
rect 1500 641 1528 1124
rect 1556 669 1584 1152
rect 1612 641 1640 1124
rect 1668 669 1696 1152
rect 1724 641 1752 1124
rect 1780 669 1808 1152
rect 1836 641 1864 1124
rect 1892 669 1920 1152
rect 1948 641 2000 1124
rect 2028 669 2056 1152
rect 2084 641 2112 1124
rect 2140 669 2168 1152
rect 2196 641 2224 1124
rect 2252 669 2280 1152
rect 2308 641 2336 1124
rect 2364 669 2392 1152
rect 2420 641 2448 1124
rect 2476 669 2504 1152
rect 2532 641 2560 1124
rect 1388 577 2560 641
rect 1388 94 1416 577
rect 1444 66 1472 549
rect 1500 94 1528 577
rect 1556 66 1584 549
rect 1612 94 1640 577
rect 1668 66 1696 549
rect 1724 94 1752 577
rect 1780 66 1808 549
rect 1836 94 1864 577
rect 1892 66 1920 549
rect 1948 94 2000 577
rect 2028 66 2056 549
rect 2084 94 2112 577
rect 2140 66 2168 549
rect 2196 94 2224 577
rect 2252 66 2280 549
rect 2308 94 2336 577
rect 2364 66 2392 549
rect 2420 94 2448 577
rect 2476 66 2504 549
rect 2532 94 2560 577
rect 2588 66 2654 1152
rect 0 0 2654 66
<< obsm2 >>
rect 0 2304 619 2370
rect 0 2220 66 2304
rect 647 2276 713 2370
rect 741 2304 1913 2370
rect 94 2248 1266 2276
rect 0 2192 619 2220
rect 0 2108 66 2192
rect 647 2164 713 2248
rect 1294 2220 1360 2304
rect 1941 2276 2007 2370
rect 2035 2304 2654 2370
rect 1388 2248 2560 2276
rect 741 2192 1913 2220
rect 94 2136 1266 2164
rect 0 2080 619 2108
rect 0 1996 66 2080
rect 647 2052 713 2136
rect 1294 2108 1360 2192
rect 1941 2164 2007 2248
rect 2588 2220 2654 2304
rect 2035 2192 2654 2220
rect 1388 2136 2560 2164
rect 741 2080 1913 2108
rect 94 2024 1266 2052
rect 0 1968 619 1996
rect 0 1884 66 1968
rect 647 1940 713 2024
rect 1294 1996 1360 2080
rect 1941 2052 2007 2136
rect 2588 2108 2654 2192
rect 2035 2080 2654 2108
rect 1388 2024 2560 2052
rect 741 1968 1913 1996
rect 94 1912 1266 1940
rect 0 1817 619 1884
rect 647 1789 713 1912
rect 1294 1884 1360 1968
rect 1941 1940 2007 2024
rect 2588 1996 2654 2080
rect 2035 1968 2654 1996
rect 1388 1912 2560 1940
rect 741 1817 1913 1884
rect 1941 1789 2007 1912
rect 2588 1884 2654 1968
rect 2035 1817 2654 1884
rect 0 1733 2654 1789
rect 0 1638 619 1705
rect 0 1554 66 1638
rect 647 1610 713 1733
rect 741 1638 1913 1705
rect 94 1582 1266 1610
rect 0 1526 619 1554
rect 0 1442 66 1526
rect 647 1498 713 1582
rect 1294 1554 1360 1638
rect 1941 1610 2007 1733
rect 2035 1638 2654 1705
rect 1388 1582 2560 1610
rect 741 1526 1913 1554
rect 94 1470 1266 1498
rect 0 1414 619 1442
rect 0 1330 66 1414
rect 647 1386 713 1470
rect 1294 1442 1360 1526
rect 1941 1498 2007 1582
rect 2588 1554 2654 1638
rect 2035 1526 2654 1554
rect 1388 1470 2560 1498
rect 741 1414 1913 1442
rect 94 1358 1266 1386
rect 0 1302 619 1330
rect 0 1218 66 1302
rect 647 1274 713 1358
rect 1294 1330 1360 1414
rect 1941 1386 2007 1470
rect 2588 1442 2654 1526
rect 2035 1414 2654 1442
rect 1388 1358 2560 1386
rect 741 1302 1913 1330
rect 94 1246 1266 1274
rect 0 1152 619 1218
rect 0 1068 66 1152
rect 647 1124 713 1246
rect 1294 1218 1360 1302
rect 1941 1274 2007 1358
rect 2588 1330 2654 1414
rect 2035 1302 2654 1330
rect 1388 1246 2560 1274
rect 741 1152 1913 1218
rect 94 1096 1266 1124
rect 0 1040 619 1068
rect 0 956 66 1040
rect 647 1012 713 1096
rect 1294 1068 1360 1152
rect 1941 1124 2007 1246
rect 2588 1218 2654 1302
rect 2035 1152 2654 1218
rect 1388 1096 2560 1124
rect 741 1040 1913 1068
rect 94 984 1266 1012
rect 0 928 619 956
rect 0 844 66 928
rect 647 900 713 984
rect 1294 956 1360 1040
rect 1941 1012 2007 1096
rect 2588 1068 2654 1152
rect 2035 1040 2654 1068
rect 1388 984 2560 1012
rect 741 928 1913 956
rect 94 872 1266 900
rect 0 816 619 844
rect 0 732 66 816
rect 647 788 713 872
rect 1294 844 1360 928
rect 1941 900 2007 984
rect 2588 956 2654 1040
rect 2035 928 2654 956
rect 1388 872 2560 900
rect 741 816 1913 844
rect 94 760 1266 788
rect 0 665 619 732
rect 647 637 713 760
rect 1294 732 1360 816
rect 1941 788 2007 872
rect 2588 844 2654 928
rect 2035 816 2654 844
rect 1388 760 2560 788
rect 741 665 1913 732
rect 1941 637 2007 760
rect 2588 732 2654 816
rect 2035 665 2654 732
rect 0 581 2654 637
rect 0 486 619 553
rect 0 402 66 486
rect 647 458 713 581
rect 741 486 1913 553
rect 94 430 1266 458
rect 0 374 619 402
rect 0 290 66 374
rect 647 346 713 430
rect 1294 402 1360 486
rect 1941 458 2007 581
rect 2035 486 2654 553
rect 1388 430 2560 458
rect 741 374 1913 402
rect 94 318 1266 346
rect 0 262 619 290
rect 0 178 66 262
rect 647 234 713 318
rect 1294 290 1360 374
rect 1941 346 2007 430
rect 2588 402 2654 486
rect 2035 374 2654 402
rect 1388 318 2560 346
rect 741 262 1913 290
rect 94 206 1266 234
rect 0 150 619 178
rect 0 66 66 150
rect 647 122 713 206
rect 1294 178 1360 262
rect 1941 234 2007 318
rect 2588 290 2654 374
rect 2035 262 2654 290
rect 1388 206 2560 234
rect 741 150 1913 178
rect 94 94 1266 122
rect 0 0 619 66
rect 647 0 713 94
rect 1294 66 1360 150
rect 1941 122 2007 206
rect 2588 178 2654 262
rect 2035 150 2654 178
rect 1388 94 2560 122
rect 741 0 1913 66
rect 1941 0 2007 94
rect 2588 66 2654 150
rect 2035 0 2654 66
<< metal3 >>
rect 0 2304 2654 2370
rect 0 1218 66 2304
rect 126 1794 194 2244
rect 254 1854 322 2304
rect 382 1794 450 2244
rect 510 1854 578 2304
rect 638 1794 722 2244
rect 782 1854 850 2304
rect 910 1794 978 2244
rect 1038 1854 1106 2304
rect 1166 1794 1234 2244
rect 126 1728 1234 1794
rect 126 1278 194 1728
rect 254 1218 322 1668
rect 382 1278 450 1728
rect 510 1218 578 1668
rect 638 1278 722 1728
rect 782 1218 850 1668
rect 910 1278 978 1728
rect 1038 1218 1106 1668
rect 1166 1278 1234 1728
rect 1294 1218 1360 2304
rect 1420 1794 1488 2244
rect 1548 1854 1616 2304
rect 1676 1794 1744 2244
rect 1804 1854 1872 2304
rect 1932 1794 2016 2244
rect 2076 1854 2144 2304
rect 2204 1794 2272 2244
rect 2332 1854 2400 2304
rect 2460 1794 2528 2244
rect 1420 1728 2528 1794
rect 1420 1278 1488 1728
rect 1548 1218 1616 1668
rect 1676 1278 1744 1728
rect 1804 1218 1872 1668
rect 1932 1278 2016 1728
rect 2076 1218 2144 1668
rect 2204 1278 2272 1728
rect 2332 1218 2400 1668
rect 2460 1278 2528 1728
rect 2588 1218 2654 2304
rect 0 1152 2654 1218
rect 0 66 66 1152
rect 126 642 194 1092
rect 254 702 322 1152
rect 382 642 450 1092
rect 510 702 578 1152
rect 638 642 722 1092
rect 782 702 850 1152
rect 910 642 978 1092
rect 1038 702 1106 1152
rect 1166 642 1234 1092
rect 126 576 1234 642
rect 126 126 194 576
rect 254 66 322 516
rect 382 126 450 576
rect 510 66 578 516
rect 638 126 722 576
rect 782 66 850 516
rect 910 126 978 576
rect 1038 66 1106 516
rect 1166 126 1234 576
rect 1294 66 1360 1152
rect 1420 642 1488 1092
rect 1548 702 1616 1152
rect 1676 642 1744 1092
rect 1804 702 1872 1152
rect 1932 642 2016 1092
rect 2076 702 2144 1152
rect 2204 642 2272 1092
rect 2332 702 2400 1152
rect 2460 642 2528 1092
rect 1420 576 2528 642
rect 1420 126 1488 576
rect 1548 66 1616 516
rect 1676 126 1744 576
rect 1804 66 1872 516
rect 1932 126 2016 576
rect 2076 66 2144 516
rect 2204 126 2272 576
rect 2332 66 2400 516
rect 2460 126 2528 576
rect 2588 66 2654 1152
rect 0 0 2654 66
<< metal4 >>
rect 0 0 2654 2370
<< labels >>
rlabel metal3 s 2588 1218 2654 2304 6 C0
port 1 nsew
rlabel metal3 s 2588 66 2654 1152 6 C0
port 1 nsew
rlabel metal3 s 2332 1854 2400 2304 6 C0
port 1 nsew
rlabel metal3 s 2332 1218 2400 1668 6 C0
port 1 nsew
rlabel metal3 s 2332 702 2400 1152 6 C0
port 1 nsew
rlabel metal3 s 2332 66 2400 516 6 C0
port 1 nsew
rlabel metal3 s 2076 1854 2144 2304 6 C0
port 1 nsew
rlabel metal3 s 2076 1218 2144 1668 6 C0
port 1 nsew
rlabel metal3 s 2076 702 2144 1152 6 C0
port 1 nsew
rlabel metal3 s 2076 66 2144 516 6 C0
port 1 nsew
rlabel metal3 s 1804 1854 1872 2304 6 C0
port 1 nsew
rlabel metal3 s 1804 1218 1872 1668 6 C0
port 1 nsew
rlabel metal3 s 1804 702 1872 1152 6 C0
port 1 nsew
rlabel metal3 s 1804 66 1872 516 6 C0
port 1 nsew
rlabel metal3 s 1548 1854 1616 2304 6 C0
port 1 nsew
rlabel metal3 s 1548 1218 1616 1668 6 C0
port 1 nsew
rlabel metal3 s 1548 702 1616 1152 6 C0
port 1 nsew
rlabel metal3 s 1548 66 1616 516 6 C0
port 1 nsew
rlabel metal3 s 1294 1218 1360 2304 6 C0
port 1 nsew
rlabel metal3 s 1294 66 1360 1152 6 C0
port 1 nsew
rlabel metal3 s 1038 1854 1106 2304 6 C0
port 1 nsew
rlabel metal3 s 1038 1218 1106 1668 6 C0
port 1 nsew
rlabel metal3 s 1038 702 1106 1152 6 C0
port 1 nsew
rlabel metal3 s 1038 66 1106 516 6 C0
port 1 nsew
rlabel metal3 s 782 1854 850 2304 6 C0
port 1 nsew
rlabel metal3 s 782 1218 850 1668 6 C0
port 1 nsew
rlabel metal3 s 782 702 850 1152 6 C0
port 1 nsew
rlabel metal3 s 782 66 850 516 6 C0
port 1 nsew
rlabel metal3 s 510 1854 578 2304 6 C0
port 1 nsew
rlabel metal3 s 510 1218 578 1668 6 C0
port 1 nsew
rlabel metal3 s 510 702 578 1152 6 C0
port 1 nsew
rlabel metal3 s 510 66 578 516 6 C0
port 1 nsew
rlabel metal3 s 254 1854 322 2304 6 C0
port 1 nsew
rlabel metal3 s 254 1218 322 1668 6 C0
port 1 nsew
rlabel metal3 s 254 702 322 1152 6 C0
port 1 nsew
rlabel metal3 s 254 66 322 516 6 C0
port 1 nsew
rlabel metal3 s 0 2304 2654 2370 6 C0
port 1 nsew
rlabel metal3 s 0 1218 66 2304 6 C0
port 1 nsew
rlabel metal3 s 0 1152 2654 1218 6 C0
port 1 nsew
rlabel metal3 s 0 66 66 1152 6 C0
port 1 nsew
rlabel metal3 s 0 0 2654 66 6 C0
port 1 nsew
rlabel metal3 s 2460 1794 2528 2244 6 C1
port 2 nsew
rlabel metal3 s 2460 1278 2528 1728 6 C1
port 2 nsew
rlabel metal3 s 2460 642 2528 1092 6 C1
port 2 nsew
rlabel metal3 s 2460 126 2528 576 6 C1
port 2 nsew
rlabel metal3 s 2204 1794 2272 2244 6 C1
port 2 nsew
rlabel metal3 s 2204 1278 2272 1728 6 C1
port 2 nsew
rlabel metal3 s 2204 642 2272 1092 6 C1
port 2 nsew
rlabel metal3 s 2204 126 2272 576 6 C1
port 2 nsew
rlabel metal3 s 1932 1794 2016 2244 6 C1
port 2 nsew
rlabel metal3 s 1932 1278 2016 1728 6 C1
port 2 nsew
rlabel metal3 s 1932 642 2016 1092 6 C1
port 2 nsew
rlabel metal3 s 1932 126 2016 576 6 C1
port 2 nsew
rlabel metal3 s 1676 1794 1744 2244 6 C1
port 2 nsew
rlabel metal3 s 1676 1278 1744 1728 6 C1
port 2 nsew
rlabel metal3 s 1676 642 1744 1092 6 C1
port 2 nsew
rlabel metal3 s 1676 126 1744 576 6 C1
port 2 nsew
rlabel metal3 s 1420 1794 1488 2244 6 C1
port 2 nsew
rlabel metal3 s 1420 1728 2528 1794 6 C1
port 2 nsew
rlabel metal3 s 1420 1278 1488 1728 6 C1
port 2 nsew
rlabel metal3 s 1420 642 1488 1092 6 C1
port 2 nsew
rlabel metal3 s 1420 576 2528 642 6 C1
port 2 nsew
rlabel metal3 s 1420 126 1488 576 6 C1
port 2 nsew
rlabel metal3 s 1166 1794 1234 2244 6 C1
port 2 nsew
rlabel metal3 s 1166 1278 1234 1728 6 C1
port 2 nsew
rlabel metal3 s 1166 642 1234 1092 6 C1
port 2 nsew
rlabel metal3 s 1166 126 1234 576 6 C1
port 2 nsew
rlabel metal3 s 910 1794 978 2244 6 C1
port 2 nsew
rlabel metal3 s 910 1278 978 1728 6 C1
port 2 nsew
rlabel metal3 s 910 642 978 1092 6 C1
port 2 nsew
rlabel metal3 s 910 126 978 576 6 C1
port 2 nsew
rlabel metal3 s 638 1794 722 2244 6 C1
port 2 nsew
rlabel metal3 s 638 1278 722 1728 6 C1
port 2 nsew
rlabel metal3 s 638 642 722 1092 6 C1
port 2 nsew
rlabel metal3 s 638 126 722 576 6 C1
port 2 nsew
rlabel metal3 s 382 1794 450 2244 6 C1
port 2 nsew
rlabel metal3 s 382 1278 450 1728 6 C1
port 2 nsew
rlabel metal3 s 382 642 450 1092 6 C1
port 2 nsew
rlabel metal3 s 382 126 450 576 6 C1
port 2 nsew
rlabel metal3 s 126 1794 194 2244 6 C1
port 2 nsew
rlabel metal3 s 126 1728 1234 1794 6 C1
port 2 nsew
rlabel metal3 s 126 1278 194 1728 6 C1
port 2 nsew
rlabel metal3 s 126 642 194 1092 6 C1
port 2 nsew
rlabel metal3 s 126 576 1234 642 6 C1
port 2 nsew
rlabel metal3 s 126 126 194 576 6 C1
port 2 nsew
rlabel metal4 s 0 0 2654 2370 6 M4
port 3 nsew
rlabel pwell s 1179 1269 1189 1279 6 SUB
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2654 2370
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 218298
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 217726
<< end >>
