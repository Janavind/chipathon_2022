magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< obsli1 >>
rect 34 2092 2158 2158
rect 34 100 100 2092
rect 260 1866 1932 1932
rect 260 326 326 1866
rect 662 1464 1530 1530
rect 662 728 728 1464
rect 893 893 1299 1299
rect 1464 728 1530 1464
rect 662 662 1530 728
rect 1866 326 1932 1866
rect 260 260 1932 326
rect 2092 100 2158 2092
rect 34 34 2158 100
<< obsm1 >>
rect 38 2096 2154 2154
rect 38 96 96 2096
rect 264 1870 1928 1928
rect 264 322 322 1870
rect 666 1468 1526 1526
rect 666 724 724 1468
rect 923 923 1269 1269
rect 1468 724 1526 1468
rect 666 666 1526 724
rect 1870 322 1928 1870
rect 264 264 1928 322
rect 2096 96 2154 2096
rect 38 38 2154 96
<< properties >>
string FIXED_BBOX 26 26 2166 2166
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8917018
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8872078
<< end >>
