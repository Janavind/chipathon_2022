magic
tech sky130B
magscale 1 2
timestamp 1666464484
use sky130_fd_pr__via_pol1__example_5595914180854  sky130_fd_pr__via_pol1__example_5595914180854_0
timestamp 1666464484
transform -1 0 16 0 1 31
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180854  sky130_fd_pr__via_pol1__example_5595914180854_1
timestamp 1666464484
transform 1 0 584 0 1 31
box 0 0 1 1
<< properties >>
string GDS_END 35992154
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 35991672
<< end >>
