magic
tech sky130B
magscale 1 2
timestamp 1666464484
use sky130_fd_pr__hvdfm1sd2__example_55959141808717  sky130_fd_pr__hvdfm1sd2__example_55959141808717_0
timestamp 1666464484
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808717  sky130_fd_pr__hvdfm1sd2__example_55959141808717_1
timestamp 1666464484
transform 1 0 200 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 3902748
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3901690
<< end >>
