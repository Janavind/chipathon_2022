magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< metal3 >>
rect 100 9930 4880 10164
rect 10151 9930 14931 10164
rect 10151 6948 14931 7636
<< obsm3 >>
rect 100 6948 4880 7636
<< metal4 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18600
rect 14746 13607 15000 18600
rect 0 12417 254 13307
rect 14746 12417 15000 13307
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 15000 10947
rect 0 10225 15000 10821
rect 0 9929 254 10165
rect 14746 9929 15000 10165
rect 0 9273 15000 9869
rect 0 9147 15000 9213
rect 0 7917 254 8847
rect 14746 7917 15000 8847
rect 0 6947 254 7637
rect 270 7568 334 7632
rect 352 7568 416 7632
rect 434 7568 498 7632
rect 516 7568 580 7632
rect 598 7568 662 7632
rect 679 7568 743 7632
rect 760 7568 824 7632
rect 841 7568 905 7632
rect 922 7568 986 7632
rect 1003 7568 1067 7632
rect 1084 7568 1148 7632
rect 1165 7568 1229 7632
rect 1246 7568 1310 7632
rect 1327 7568 1391 7632
rect 1408 7568 1472 7632
rect 1489 7568 1553 7632
rect 1570 7568 1634 7632
rect 1651 7568 1715 7632
rect 1732 7568 1796 7632
rect 1813 7568 1877 7632
rect 1894 7568 1958 7632
rect 1975 7568 2039 7632
rect 2056 7568 2120 7632
rect 2137 7568 2201 7632
rect 2218 7568 2282 7632
rect 2299 7568 2363 7632
rect 2380 7568 2444 7632
rect 2461 7568 2525 7632
rect 2542 7568 2606 7632
rect 2623 7568 2687 7632
rect 2704 7568 2768 7632
rect 2785 7568 2849 7632
rect 2866 7568 2930 7632
rect 2947 7568 3011 7632
rect 3028 7568 3092 7632
rect 3109 7568 3173 7632
rect 3190 7568 3254 7632
rect 3271 7568 3335 7632
rect 3352 7568 3416 7632
rect 3433 7568 3497 7632
rect 3514 7568 3578 7632
rect 3595 7568 3659 7632
rect 3676 7568 3740 7632
rect 3757 7568 3821 7632
rect 3838 7568 3902 7632
rect 3919 7568 3983 7632
rect 4000 7568 4064 7632
rect 4081 7568 4145 7632
rect 4162 7568 4226 7632
rect 4243 7568 4307 7632
rect 4324 7568 4388 7632
rect 4405 7568 4469 7632
rect 4486 7568 4550 7632
rect 4567 7568 4631 7632
rect 4648 7568 4712 7632
rect 4729 7568 4793 7632
rect 4810 7568 4874 7632
rect 270 7480 334 7544
rect 352 7480 416 7544
rect 434 7480 498 7544
rect 516 7480 580 7544
rect 598 7480 662 7544
rect 679 7480 743 7544
rect 760 7480 824 7544
rect 841 7480 905 7544
rect 922 7480 986 7544
rect 1003 7480 1067 7544
rect 1084 7480 1148 7544
rect 1165 7480 1229 7544
rect 1246 7480 1310 7544
rect 1327 7480 1391 7544
rect 1408 7480 1472 7544
rect 1489 7480 1553 7544
rect 1570 7480 1634 7544
rect 1651 7480 1715 7544
rect 1732 7480 1796 7544
rect 1813 7480 1877 7544
rect 1894 7480 1958 7544
rect 1975 7480 2039 7544
rect 2056 7480 2120 7544
rect 2137 7480 2201 7544
rect 2218 7480 2282 7544
rect 2299 7480 2363 7544
rect 2380 7480 2444 7544
rect 2461 7480 2525 7544
rect 2542 7480 2606 7544
rect 2623 7480 2687 7544
rect 2704 7480 2768 7544
rect 2785 7480 2849 7544
rect 2866 7480 2930 7544
rect 2947 7480 3011 7544
rect 3028 7480 3092 7544
rect 3109 7480 3173 7544
rect 3190 7480 3254 7544
rect 3271 7480 3335 7544
rect 3352 7480 3416 7544
rect 3433 7480 3497 7544
rect 3514 7480 3578 7544
rect 3595 7480 3659 7544
rect 3676 7480 3740 7544
rect 3757 7480 3821 7544
rect 3838 7480 3902 7544
rect 3919 7480 3983 7544
rect 4000 7480 4064 7544
rect 4081 7480 4145 7544
rect 4162 7480 4226 7544
rect 4243 7480 4307 7544
rect 4324 7480 4388 7544
rect 4405 7480 4469 7544
rect 4486 7480 4550 7544
rect 4567 7480 4631 7544
rect 4648 7480 4712 7544
rect 4729 7480 4793 7544
rect 4810 7480 4874 7544
rect 270 7392 334 7456
rect 352 7392 416 7456
rect 434 7392 498 7456
rect 516 7392 580 7456
rect 598 7392 662 7456
rect 679 7392 743 7456
rect 760 7392 824 7456
rect 841 7392 905 7456
rect 922 7392 986 7456
rect 1003 7392 1067 7456
rect 1084 7392 1148 7456
rect 1165 7392 1229 7456
rect 1246 7392 1310 7456
rect 1327 7392 1391 7456
rect 1408 7392 1472 7456
rect 1489 7392 1553 7456
rect 1570 7392 1634 7456
rect 1651 7392 1715 7456
rect 1732 7392 1796 7456
rect 1813 7392 1877 7456
rect 1894 7392 1958 7456
rect 1975 7392 2039 7456
rect 2056 7392 2120 7456
rect 2137 7392 2201 7456
rect 2218 7392 2282 7456
rect 2299 7392 2363 7456
rect 2380 7392 2444 7456
rect 2461 7392 2525 7456
rect 2542 7392 2606 7456
rect 2623 7392 2687 7456
rect 2704 7392 2768 7456
rect 2785 7392 2849 7456
rect 2866 7392 2930 7456
rect 2947 7392 3011 7456
rect 3028 7392 3092 7456
rect 3109 7392 3173 7456
rect 3190 7392 3254 7456
rect 3271 7392 3335 7456
rect 3352 7392 3416 7456
rect 3433 7392 3497 7456
rect 3514 7392 3578 7456
rect 3595 7392 3659 7456
rect 3676 7392 3740 7456
rect 3757 7392 3821 7456
rect 3838 7392 3902 7456
rect 3919 7392 3983 7456
rect 4000 7392 4064 7456
rect 4081 7392 4145 7456
rect 4162 7392 4226 7456
rect 4243 7392 4307 7456
rect 4324 7392 4388 7456
rect 4405 7392 4469 7456
rect 4486 7392 4550 7456
rect 4567 7392 4631 7456
rect 4648 7392 4712 7456
rect 4729 7392 4793 7456
rect 4810 7392 4874 7456
rect 270 7304 334 7368
rect 352 7304 416 7368
rect 434 7304 498 7368
rect 516 7304 580 7368
rect 598 7304 662 7368
rect 679 7304 743 7368
rect 760 7304 824 7368
rect 841 7304 905 7368
rect 922 7304 986 7368
rect 1003 7304 1067 7368
rect 1084 7304 1148 7368
rect 1165 7304 1229 7368
rect 1246 7304 1310 7368
rect 1327 7304 1391 7368
rect 1408 7304 1472 7368
rect 1489 7304 1553 7368
rect 1570 7304 1634 7368
rect 1651 7304 1715 7368
rect 1732 7304 1796 7368
rect 1813 7304 1877 7368
rect 1894 7304 1958 7368
rect 1975 7304 2039 7368
rect 2056 7304 2120 7368
rect 2137 7304 2201 7368
rect 2218 7304 2282 7368
rect 2299 7304 2363 7368
rect 2380 7304 2444 7368
rect 2461 7304 2525 7368
rect 2542 7304 2606 7368
rect 2623 7304 2687 7368
rect 2704 7304 2768 7368
rect 2785 7304 2849 7368
rect 2866 7304 2930 7368
rect 2947 7304 3011 7368
rect 3028 7304 3092 7368
rect 3109 7304 3173 7368
rect 3190 7304 3254 7368
rect 3271 7304 3335 7368
rect 3352 7304 3416 7368
rect 3433 7304 3497 7368
rect 3514 7304 3578 7368
rect 3595 7304 3659 7368
rect 3676 7304 3740 7368
rect 3757 7304 3821 7368
rect 3838 7304 3902 7368
rect 3919 7304 3983 7368
rect 4000 7304 4064 7368
rect 4081 7304 4145 7368
rect 4162 7304 4226 7368
rect 4243 7304 4307 7368
rect 4324 7304 4388 7368
rect 4405 7304 4469 7368
rect 4486 7304 4550 7368
rect 4567 7304 4631 7368
rect 4648 7304 4712 7368
rect 4729 7304 4793 7368
rect 4810 7304 4874 7368
rect 270 7216 334 7280
rect 352 7216 416 7280
rect 434 7216 498 7280
rect 516 7216 580 7280
rect 598 7216 662 7280
rect 679 7216 743 7280
rect 760 7216 824 7280
rect 841 7216 905 7280
rect 922 7216 986 7280
rect 1003 7216 1067 7280
rect 1084 7216 1148 7280
rect 1165 7216 1229 7280
rect 1246 7216 1310 7280
rect 1327 7216 1391 7280
rect 1408 7216 1472 7280
rect 1489 7216 1553 7280
rect 1570 7216 1634 7280
rect 1651 7216 1715 7280
rect 1732 7216 1796 7280
rect 1813 7216 1877 7280
rect 1894 7216 1958 7280
rect 1975 7216 2039 7280
rect 2056 7216 2120 7280
rect 2137 7216 2201 7280
rect 2218 7216 2282 7280
rect 2299 7216 2363 7280
rect 2380 7216 2444 7280
rect 2461 7216 2525 7280
rect 2542 7216 2606 7280
rect 2623 7216 2687 7280
rect 2704 7216 2768 7280
rect 2785 7216 2849 7280
rect 2866 7216 2930 7280
rect 2947 7216 3011 7280
rect 3028 7216 3092 7280
rect 3109 7216 3173 7280
rect 3190 7216 3254 7280
rect 3271 7216 3335 7280
rect 3352 7216 3416 7280
rect 3433 7216 3497 7280
rect 3514 7216 3578 7280
rect 3595 7216 3659 7280
rect 3676 7216 3740 7280
rect 3757 7216 3821 7280
rect 3838 7216 3902 7280
rect 3919 7216 3983 7280
rect 4000 7216 4064 7280
rect 4081 7216 4145 7280
rect 4162 7216 4226 7280
rect 4243 7216 4307 7280
rect 4324 7216 4388 7280
rect 4405 7216 4469 7280
rect 4486 7216 4550 7280
rect 4567 7216 4631 7280
rect 4648 7216 4712 7280
rect 4729 7216 4793 7280
rect 4810 7216 4874 7280
rect 270 7128 334 7192
rect 352 7128 416 7192
rect 434 7128 498 7192
rect 516 7128 580 7192
rect 598 7128 662 7192
rect 679 7128 743 7192
rect 760 7128 824 7192
rect 841 7128 905 7192
rect 922 7128 986 7192
rect 1003 7128 1067 7192
rect 1084 7128 1148 7192
rect 1165 7128 1229 7192
rect 1246 7128 1310 7192
rect 1327 7128 1391 7192
rect 1408 7128 1472 7192
rect 1489 7128 1553 7192
rect 1570 7128 1634 7192
rect 1651 7128 1715 7192
rect 1732 7128 1796 7192
rect 1813 7128 1877 7192
rect 1894 7128 1958 7192
rect 1975 7128 2039 7192
rect 2056 7128 2120 7192
rect 2137 7128 2201 7192
rect 2218 7128 2282 7192
rect 2299 7128 2363 7192
rect 2380 7128 2444 7192
rect 2461 7128 2525 7192
rect 2542 7128 2606 7192
rect 2623 7128 2687 7192
rect 2704 7128 2768 7192
rect 2785 7128 2849 7192
rect 2866 7128 2930 7192
rect 2947 7128 3011 7192
rect 3028 7128 3092 7192
rect 3109 7128 3173 7192
rect 3190 7128 3254 7192
rect 3271 7128 3335 7192
rect 3352 7128 3416 7192
rect 3433 7128 3497 7192
rect 3514 7128 3578 7192
rect 3595 7128 3659 7192
rect 3676 7128 3740 7192
rect 3757 7128 3821 7192
rect 3838 7128 3902 7192
rect 3919 7128 3983 7192
rect 4000 7128 4064 7192
rect 4081 7128 4145 7192
rect 4162 7128 4226 7192
rect 4243 7128 4307 7192
rect 4324 7128 4388 7192
rect 4405 7128 4469 7192
rect 4486 7128 4550 7192
rect 4567 7128 4631 7192
rect 4648 7128 4712 7192
rect 4729 7128 4793 7192
rect 4810 7128 4874 7192
rect 270 7040 334 7104
rect 352 7040 416 7104
rect 434 7040 498 7104
rect 516 7040 580 7104
rect 598 7040 662 7104
rect 679 7040 743 7104
rect 760 7040 824 7104
rect 841 7040 905 7104
rect 922 7040 986 7104
rect 1003 7040 1067 7104
rect 1084 7040 1148 7104
rect 1165 7040 1229 7104
rect 1246 7040 1310 7104
rect 1327 7040 1391 7104
rect 1408 7040 1472 7104
rect 1489 7040 1553 7104
rect 1570 7040 1634 7104
rect 1651 7040 1715 7104
rect 1732 7040 1796 7104
rect 1813 7040 1877 7104
rect 1894 7040 1958 7104
rect 1975 7040 2039 7104
rect 2056 7040 2120 7104
rect 2137 7040 2201 7104
rect 2218 7040 2282 7104
rect 2299 7040 2363 7104
rect 2380 7040 2444 7104
rect 2461 7040 2525 7104
rect 2542 7040 2606 7104
rect 2623 7040 2687 7104
rect 2704 7040 2768 7104
rect 2785 7040 2849 7104
rect 2866 7040 2930 7104
rect 2947 7040 3011 7104
rect 3028 7040 3092 7104
rect 3109 7040 3173 7104
rect 3190 7040 3254 7104
rect 3271 7040 3335 7104
rect 3352 7040 3416 7104
rect 3433 7040 3497 7104
rect 3514 7040 3578 7104
rect 3595 7040 3659 7104
rect 3676 7040 3740 7104
rect 3757 7040 3821 7104
rect 3838 7040 3902 7104
rect 3919 7040 3983 7104
rect 4000 7040 4064 7104
rect 4081 7040 4145 7104
rect 4162 7040 4226 7104
rect 4243 7040 4307 7104
rect 4324 7040 4388 7104
rect 4405 7040 4469 7104
rect 4486 7040 4550 7104
rect 4567 7040 4631 7104
rect 4648 7040 4712 7104
rect 4729 7040 4793 7104
rect 4810 7040 4874 7104
rect 270 6952 334 7016
rect 352 6952 416 7016
rect 434 6952 498 7016
rect 516 6952 580 7016
rect 598 6952 662 7016
rect 679 6952 743 7016
rect 760 6952 824 7016
rect 841 6952 905 7016
rect 922 6952 986 7016
rect 1003 6952 1067 7016
rect 1084 6952 1148 7016
rect 1165 6952 1229 7016
rect 1246 6952 1310 7016
rect 1327 6952 1391 7016
rect 1408 6952 1472 7016
rect 1489 6952 1553 7016
rect 1570 6952 1634 7016
rect 1651 6952 1715 7016
rect 1732 6952 1796 7016
rect 1813 6952 1877 7016
rect 1894 6952 1958 7016
rect 1975 6952 2039 7016
rect 2056 6952 2120 7016
rect 2137 6952 2201 7016
rect 2218 6952 2282 7016
rect 2299 6952 2363 7016
rect 2380 6952 2444 7016
rect 2461 6952 2525 7016
rect 2542 6952 2606 7016
rect 2623 6952 2687 7016
rect 2704 6952 2768 7016
rect 2785 6952 2849 7016
rect 2866 6952 2930 7016
rect 2947 6952 3011 7016
rect 3028 6952 3092 7016
rect 3109 6952 3173 7016
rect 3190 6952 3254 7016
rect 3271 6952 3335 7016
rect 3352 6952 3416 7016
rect 3433 6952 3497 7016
rect 3514 6952 3578 7016
rect 3595 6952 3659 7016
rect 3676 6952 3740 7016
rect 3757 6952 3821 7016
rect 3838 6952 3902 7016
rect 3919 6952 3983 7016
rect 4000 6952 4064 7016
rect 4081 6952 4145 7016
rect 4162 6952 4226 7016
rect 4243 6952 4307 7016
rect 4324 6952 4388 7016
rect 4405 6952 4469 7016
rect 4486 6952 4550 7016
rect 4567 6952 4631 7016
rect 4648 6952 4712 7016
rect 4729 6952 4793 7016
rect 4810 6952 4874 7016
rect 14746 6947 15000 7637
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 14746 4767 15000 5697
rect 0 3557 254 4487
rect 14746 3557 15000 4487
rect 0 2587 193 3277
rect 14807 2587 15000 3277
rect 0 1377 254 2307
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< obsm4 >>
rect 334 34677 14666 39600
rect 193 18680 14807 34677
rect 334 13527 14666 18680
rect 193 13387 14807 13527
rect 334 12337 14666 13387
rect 193 12217 14807 12337
rect 334 11167 14666 12217
rect 193 11027 14807 11167
rect 334 9949 14666 10145
rect 193 8927 14807 9067
rect 334 7837 14666 8927
rect 193 7717 14807 7837
rect 334 7632 14666 7717
rect 334 7568 352 7632
rect 416 7568 434 7632
rect 498 7568 516 7632
rect 580 7568 598 7632
rect 662 7568 679 7632
rect 743 7568 760 7632
rect 824 7568 841 7632
rect 905 7568 922 7632
rect 986 7568 1003 7632
rect 1067 7568 1084 7632
rect 1148 7568 1165 7632
rect 1229 7568 1246 7632
rect 1310 7568 1327 7632
rect 1391 7568 1408 7632
rect 1472 7568 1489 7632
rect 1553 7568 1570 7632
rect 1634 7568 1651 7632
rect 1715 7568 1732 7632
rect 1796 7568 1813 7632
rect 1877 7568 1894 7632
rect 1958 7568 1975 7632
rect 2039 7568 2056 7632
rect 2120 7568 2137 7632
rect 2201 7568 2218 7632
rect 2282 7568 2299 7632
rect 2363 7568 2380 7632
rect 2444 7568 2461 7632
rect 2525 7568 2542 7632
rect 2606 7568 2623 7632
rect 2687 7568 2704 7632
rect 2768 7568 2785 7632
rect 2849 7568 2866 7632
rect 2930 7568 2947 7632
rect 3011 7568 3028 7632
rect 3092 7568 3109 7632
rect 3173 7568 3190 7632
rect 3254 7568 3271 7632
rect 3335 7568 3352 7632
rect 3416 7568 3433 7632
rect 3497 7568 3514 7632
rect 3578 7568 3595 7632
rect 3659 7568 3676 7632
rect 3740 7568 3757 7632
rect 3821 7568 3838 7632
rect 3902 7568 3919 7632
rect 3983 7568 4000 7632
rect 4064 7568 4081 7632
rect 4145 7568 4162 7632
rect 4226 7568 4243 7632
rect 4307 7568 4324 7632
rect 4388 7568 4405 7632
rect 4469 7568 4486 7632
rect 4550 7568 4567 7632
rect 4631 7568 4648 7632
rect 4712 7568 4729 7632
rect 4793 7568 4810 7632
rect 4874 7568 14666 7632
rect 334 7544 14666 7568
rect 334 7480 352 7544
rect 416 7480 434 7544
rect 498 7480 516 7544
rect 580 7480 598 7544
rect 662 7480 679 7544
rect 743 7480 760 7544
rect 824 7480 841 7544
rect 905 7480 922 7544
rect 986 7480 1003 7544
rect 1067 7480 1084 7544
rect 1148 7480 1165 7544
rect 1229 7480 1246 7544
rect 1310 7480 1327 7544
rect 1391 7480 1408 7544
rect 1472 7480 1489 7544
rect 1553 7480 1570 7544
rect 1634 7480 1651 7544
rect 1715 7480 1732 7544
rect 1796 7480 1813 7544
rect 1877 7480 1894 7544
rect 1958 7480 1975 7544
rect 2039 7480 2056 7544
rect 2120 7480 2137 7544
rect 2201 7480 2218 7544
rect 2282 7480 2299 7544
rect 2363 7480 2380 7544
rect 2444 7480 2461 7544
rect 2525 7480 2542 7544
rect 2606 7480 2623 7544
rect 2687 7480 2704 7544
rect 2768 7480 2785 7544
rect 2849 7480 2866 7544
rect 2930 7480 2947 7544
rect 3011 7480 3028 7544
rect 3092 7480 3109 7544
rect 3173 7480 3190 7544
rect 3254 7480 3271 7544
rect 3335 7480 3352 7544
rect 3416 7480 3433 7544
rect 3497 7480 3514 7544
rect 3578 7480 3595 7544
rect 3659 7480 3676 7544
rect 3740 7480 3757 7544
rect 3821 7480 3838 7544
rect 3902 7480 3919 7544
rect 3983 7480 4000 7544
rect 4064 7480 4081 7544
rect 4145 7480 4162 7544
rect 4226 7480 4243 7544
rect 4307 7480 4324 7544
rect 4388 7480 4405 7544
rect 4469 7480 4486 7544
rect 4550 7480 4567 7544
rect 4631 7480 4648 7544
rect 4712 7480 4729 7544
rect 4793 7480 4810 7544
rect 4874 7480 14666 7544
rect 334 7456 14666 7480
rect 334 7392 352 7456
rect 416 7392 434 7456
rect 498 7392 516 7456
rect 580 7392 598 7456
rect 662 7392 679 7456
rect 743 7392 760 7456
rect 824 7392 841 7456
rect 905 7392 922 7456
rect 986 7392 1003 7456
rect 1067 7392 1084 7456
rect 1148 7392 1165 7456
rect 1229 7392 1246 7456
rect 1310 7392 1327 7456
rect 1391 7392 1408 7456
rect 1472 7392 1489 7456
rect 1553 7392 1570 7456
rect 1634 7392 1651 7456
rect 1715 7392 1732 7456
rect 1796 7392 1813 7456
rect 1877 7392 1894 7456
rect 1958 7392 1975 7456
rect 2039 7392 2056 7456
rect 2120 7392 2137 7456
rect 2201 7392 2218 7456
rect 2282 7392 2299 7456
rect 2363 7392 2380 7456
rect 2444 7392 2461 7456
rect 2525 7392 2542 7456
rect 2606 7392 2623 7456
rect 2687 7392 2704 7456
rect 2768 7392 2785 7456
rect 2849 7392 2866 7456
rect 2930 7392 2947 7456
rect 3011 7392 3028 7456
rect 3092 7392 3109 7456
rect 3173 7392 3190 7456
rect 3254 7392 3271 7456
rect 3335 7392 3352 7456
rect 3416 7392 3433 7456
rect 3497 7392 3514 7456
rect 3578 7392 3595 7456
rect 3659 7392 3676 7456
rect 3740 7392 3757 7456
rect 3821 7392 3838 7456
rect 3902 7392 3919 7456
rect 3983 7392 4000 7456
rect 4064 7392 4081 7456
rect 4145 7392 4162 7456
rect 4226 7392 4243 7456
rect 4307 7392 4324 7456
rect 4388 7392 4405 7456
rect 4469 7392 4486 7456
rect 4550 7392 4567 7456
rect 4631 7392 4648 7456
rect 4712 7392 4729 7456
rect 4793 7392 4810 7456
rect 4874 7392 14666 7456
rect 334 7368 14666 7392
rect 334 7304 352 7368
rect 416 7304 434 7368
rect 498 7304 516 7368
rect 580 7304 598 7368
rect 662 7304 679 7368
rect 743 7304 760 7368
rect 824 7304 841 7368
rect 905 7304 922 7368
rect 986 7304 1003 7368
rect 1067 7304 1084 7368
rect 1148 7304 1165 7368
rect 1229 7304 1246 7368
rect 1310 7304 1327 7368
rect 1391 7304 1408 7368
rect 1472 7304 1489 7368
rect 1553 7304 1570 7368
rect 1634 7304 1651 7368
rect 1715 7304 1732 7368
rect 1796 7304 1813 7368
rect 1877 7304 1894 7368
rect 1958 7304 1975 7368
rect 2039 7304 2056 7368
rect 2120 7304 2137 7368
rect 2201 7304 2218 7368
rect 2282 7304 2299 7368
rect 2363 7304 2380 7368
rect 2444 7304 2461 7368
rect 2525 7304 2542 7368
rect 2606 7304 2623 7368
rect 2687 7304 2704 7368
rect 2768 7304 2785 7368
rect 2849 7304 2866 7368
rect 2930 7304 2947 7368
rect 3011 7304 3028 7368
rect 3092 7304 3109 7368
rect 3173 7304 3190 7368
rect 3254 7304 3271 7368
rect 3335 7304 3352 7368
rect 3416 7304 3433 7368
rect 3497 7304 3514 7368
rect 3578 7304 3595 7368
rect 3659 7304 3676 7368
rect 3740 7304 3757 7368
rect 3821 7304 3838 7368
rect 3902 7304 3919 7368
rect 3983 7304 4000 7368
rect 4064 7304 4081 7368
rect 4145 7304 4162 7368
rect 4226 7304 4243 7368
rect 4307 7304 4324 7368
rect 4388 7304 4405 7368
rect 4469 7304 4486 7368
rect 4550 7304 4567 7368
rect 4631 7304 4648 7368
rect 4712 7304 4729 7368
rect 4793 7304 4810 7368
rect 4874 7304 14666 7368
rect 334 7280 14666 7304
rect 334 7216 352 7280
rect 416 7216 434 7280
rect 498 7216 516 7280
rect 580 7216 598 7280
rect 662 7216 679 7280
rect 743 7216 760 7280
rect 824 7216 841 7280
rect 905 7216 922 7280
rect 986 7216 1003 7280
rect 1067 7216 1084 7280
rect 1148 7216 1165 7280
rect 1229 7216 1246 7280
rect 1310 7216 1327 7280
rect 1391 7216 1408 7280
rect 1472 7216 1489 7280
rect 1553 7216 1570 7280
rect 1634 7216 1651 7280
rect 1715 7216 1732 7280
rect 1796 7216 1813 7280
rect 1877 7216 1894 7280
rect 1958 7216 1975 7280
rect 2039 7216 2056 7280
rect 2120 7216 2137 7280
rect 2201 7216 2218 7280
rect 2282 7216 2299 7280
rect 2363 7216 2380 7280
rect 2444 7216 2461 7280
rect 2525 7216 2542 7280
rect 2606 7216 2623 7280
rect 2687 7216 2704 7280
rect 2768 7216 2785 7280
rect 2849 7216 2866 7280
rect 2930 7216 2947 7280
rect 3011 7216 3028 7280
rect 3092 7216 3109 7280
rect 3173 7216 3190 7280
rect 3254 7216 3271 7280
rect 3335 7216 3352 7280
rect 3416 7216 3433 7280
rect 3497 7216 3514 7280
rect 3578 7216 3595 7280
rect 3659 7216 3676 7280
rect 3740 7216 3757 7280
rect 3821 7216 3838 7280
rect 3902 7216 3919 7280
rect 3983 7216 4000 7280
rect 4064 7216 4081 7280
rect 4145 7216 4162 7280
rect 4226 7216 4243 7280
rect 4307 7216 4324 7280
rect 4388 7216 4405 7280
rect 4469 7216 4486 7280
rect 4550 7216 4567 7280
rect 4631 7216 4648 7280
rect 4712 7216 4729 7280
rect 4793 7216 4810 7280
rect 4874 7216 14666 7280
rect 334 7192 14666 7216
rect 334 7128 352 7192
rect 416 7128 434 7192
rect 498 7128 516 7192
rect 580 7128 598 7192
rect 662 7128 679 7192
rect 743 7128 760 7192
rect 824 7128 841 7192
rect 905 7128 922 7192
rect 986 7128 1003 7192
rect 1067 7128 1084 7192
rect 1148 7128 1165 7192
rect 1229 7128 1246 7192
rect 1310 7128 1327 7192
rect 1391 7128 1408 7192
rect 1472 7128 1489 7192
rect 1553 7128 1570 7192
rect 1634 7128 1651 7192
rect 1715 7128 1732 7192
rect 1796 7128 1813 7192
rect 1877 7128 1894 7192
rect 1958 7128 1975 7192
rect 2039 7128 2056 7192
rect 2120 7128 2137 7192
rect 2201 7128 2218 7192
rect 2282 7128 2299 7192
rect 2363 7128 2380 7192
rect 2444 7128 2461 7192
rect 2525 7128 2542 7192
rect 2606 7128 2623 7192
rect 2687 7128 2704 7192
rect 2768 7128 2785 7192
rect 2849 7128 2866 7192
rect 2930 7128 2947 7192
rect 3011 7128 3028 7192
rect 3092 7128 3109 7192
rect 3173 7128 3190 7192
rect 3254 7128 3271 7192
rect 3335 7128 3352 7192
rect 3416 7128 3433 7192
rect 3497 7128 3514 7192
rect 3578 7128 3595 7192
rect 3659 7128 3676 7192
rect 3740 7128 3757 7192
rect 3821 7128 3838 7192
rect 3902 7128 3919 7192
rect 3983 7128 4000 7192
rect 4064 7128 4081 7192
rect 4145 7128 4162 7192
rect 4226 7128 4243 7192
rect 4307 7128 4324 7192
rect 4388 7128 4405 7192
rect 4469 7128 4486 7192
rect 4550 7128 4567 7192
rect 4631 7128 4648 7192
rect 4712 7128 4729 7192
rect 4793 7128 4810 7192
rect 4874 7128 14666 7192
rect 334 7104 14666 7128
rect 334 7040 352 7104
rect 416 7040 434 7104
rect 498 7040 516 7104
rect 580 7040 598 7104
rect 662 7040 679 7104
rect 743 7040 760 7104
rect 824 7040 841 7104
rect 905 7040 922 7104
rect 986 7040 1003 7104
rect 1067 7040 1084 7104
rect 1148 7040 1165 7104
rect 1229 7040 1246 7104
rect 1310 7040 1327 7104
rect 1391 7040 1408 7104
rect 1472 7040 1489 7104
rect 1553 7040 1570 7104
rect 1634 7040 1651 7104
rect 1715 7040 1732 7104
rect 1796 7040 1813 7104
rect 1877 7040 1894 7104
rect 1958 7040 1975 7104
rect 2039 7040 2056 7104
rect 2120 7040 2137 7104
rect 2201 7040 2218 7104
rect 2282 7040 2299 7104
rect 2363 7040 2380 7104
rect 2444 7040 2461 7104
rect 2525 7040 2542 7104
rect 2606 7040 2623 7104
rect 2687 7040 2704 7104
rect 2768 7040 2785 7104
rect 2849 7040 2866 7104
rect 2930 7040 2947 7104
rect 3011 7040 3028 7104
rect 3092 7040 3109 7104
rect 3173 7040 3190 7104
rect 3254 7040 3271 7104
rect 3335 7040 3352 7104
rect 3416 7040 3433 7104
rect 3497 7040 3514 7104
rect 3578 7040 3595 7104
rect 3659 7040 3676 7104
rect 3740 7040 3757 7104
rect 3821 7040 3838 7104
rect 3902 7040 3919 7104
rect 3983 7040 4000 7104
rect 4064 7040 4081 7104
rect 4145 7040 4162 7104
rect 4226 7040 4243 7104
rect 4307 7040 4324 7104
rect 4388 7040 4405 7104
rect 4469 7040 4486 7104
rect 4550 7040 4567 7104
rect 4631 7040 4648 7104
rect 4712 7040 4729 7104
rect 4793 7040 4810 7104
rect 4874 7040 14666 7104
rect 334 7016 14666 7040
rect 334 6952 352 7016
rect 416 6952 434 7016
rect 498 6952 516 7016
rect 580 6952 598 7016
rect 662 6952 679 7016
rect 743 6952 760 7016
rect 824 6952 841 7016
rect 905 6952 922 7016
rect 986 6952 1003 7016
rect 1067 6952 1084 7016
rect 1148 6952 1165 7016
rect 1229 6952 1246 7016
rect 1310 6952 1327 7016
rect 1391 6952 1408 7016
rect 1472 6952 1489 7016
rect 1553 6952 1570 7016
rect 1634 6952 1651 7016
rect 1715 6952 1732 7016
rect 1796 6952 1813 7016
rect 1877 6952 1894 7016
rect 1958 6952 1975 7016
rect 2039 6952 2056 7016
rect 2120 6952 2137 7016
rect 2201 6952 2218 7016
rect 2282 6952 2299 7016
rect 2363 6952 2380 7016
rect 2444 6952 2461 7016
rect 2525 6952 2542 7016
rect 2606 6952 2623 7016
rect 2687 6952 2704 7016
rect 2768 6952 2785 7016
rect 2849 6952 2866 7016
rect 2930 6952 2947 7016
rect 3011 6952 3028 7016
rect 3092 6952 3109 7016
rect 3173 6952 3190 7016
rect 3254 6952 3271 7016
rect 3335 6952 3352 7016
rect 3416 6952 3433 7016
rect 3497 6952 3514 7016
rect 3578 6952 3595 7016
rect 3659 6952 3676 7016
rect 3740 6952 3757 7016
rect 3821 6952 3838 7016
rect 3902 6952 3919 7016
rect 3983 6952 4000 7016
rect 4064 6952 4081 7016
rect 4145 6952 4162 7016
rect 4226 6952 4243 7016
rect 4307 6952 4324 7016
rect 4388 6952 4405 7016
rect 4469 6952 4486 7016
rect 4550 6952 4567 7016
rect 4631 6952 4648 7016
rect 4712 6952 4729 7016
rect 4793 6952 4810 7016
rect 4874 6952 14666 7016
rect 334 6867 14666 6952
rect 193 6747 14807 6867
rect 334 5897 14666 6747
rect 193 5777 14807 5897
rect 334 4687 14666 5777
rect 193 4567 14807 4687
rect 334 3477 14666 4567
rect 193 3357 14807 3477
rect 273 2507 14727 3357
rect 193 2387 14807 2507
rect 334 1297 14666 2387
rect 193 1177 14807 1297
rect 334 7 14666 1177
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18597
rect 0 12437 254 13287
rect 0 11267 254 12117
rect 0 9147 254 10947
rect 0 7937 254 8827
rect 0 6968 254 7617
rect 14746 13607 15000 18597
rect 14746 12437 15000 13287
rect 14746 11267 15000 12117
rect 14746 9147 15000 10947
rect 14746 7937 15000 8827
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 0 4787 254 5677
rect 0 3577 254 4467
rect 14746 5997 15000 6647
rect 14746 4787 15000 5677
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 0 27 254 1077
rect 14746 1397 15000 2287
rect 14746 27 15000 1077
<< obsm5 >>
rect 574 34437 14426 39600
rect 0 18917 15000 34437
rect 574 6968 14426 18917
rect 0 6967 15000 6968
rect 574 3257 14426 6967
rect 513 2607 14487 3257
rect 574 27 14426 2607
<< labels >>
rlabel metal5 s 0 12437 254 13287 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 0 12417 254 13307 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 VSSA
port 2 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 6 VSSA
port 2 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 6 VSSA
port 2 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 0 9147 15000 9213 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 0 10881 15000 10947 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 0 6947 254 7637 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 100 9930 4880 10164 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10151 6948 14931 7636 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10151 9930 14931 10164 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14873 10111 14913 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14873 10027 14913 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14873 9943 14913 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14873 7580 14913 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14873 7492 14913 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14873 7404 14913 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14873 7316 14913 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14873 7228 14913 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14873 7140 14913 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14873 7052 14913 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14873 6964 14913 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14792 10111 14832 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14792 10027 14832 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14792 9943 14832 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14792 7580 14832 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14792 7492 14832 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14792 7404 14832 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14792 7316 14832 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14792 7228 14832 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14792 7140 14832 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14792 7052 14832 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14792 6964 14832 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14711 10111 14751 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14711 10027 14751 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14711 9943 14751 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14711 7580 14751 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14711 7492 14751 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14711 7404 14751 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14711 7316 14751 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14711 7228 14751 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14711 7140 14751 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14711 7052 14751 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14711 6964 14751 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14630 10111 14670 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14630 10027 14670 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14630 9943 14670 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14630 7580 14670 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14630 7492 14670 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14630 7404 14670 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14630 7316 14670 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14630 7228 14670 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14630 7140 14670 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14630 7052 14670 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14630 6964 14670 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14549 10111 14589 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14549 10027 14589 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14549 9943 14589 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14549 7580 14589 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14549 7492 14589 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14549 7404 14589 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14549 7316 14589 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14549 7228 14589 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14549 7140 14589 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14549 7052 14589 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14549 6964 14589 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14468 10111 14508 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14468 10027 14508 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14468 9943 14508 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14468 7580 14508 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14468 7492 14508 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14468 7404 14508 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14468 7316 14508 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14468 7228 14508 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14468 7140 14508 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14468 7052 14508 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14468 6964 14508 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14387 10111 14427 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14387 10027 14427 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14387 9943 14427 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14387 7580 14427 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14387 7492 14427 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14387 7404 14427 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14387 7316 14427 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14387 7228 14427 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14387 7140 14427 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14387 7052 14427 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14387 6964 14427 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14306 10111 14346 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14306 10027 14346 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14306 9943 14346 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14306 7580 14346 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14306 7492 14346 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14306 7404 14346 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14306 7316 14346 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14306 7228 14346 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14306 7140 14346 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14306 7052 14346 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14306 6964 14346 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14225 10111 14265 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14225 10027 14265 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14225 9943 14265 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14225 7580 14265 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14225 7492 14265 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14225 7404 14265 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14225 7316 14265 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14225 7228 14265 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14225 7140 14265 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14225 7052 14265 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14225 6964 14265 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14144 10111 14184 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14144 10027 14184 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14144 9943 14184 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14144 7580 14184 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14144 7492 14184 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14144 7404 14184 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14144 7316 14184 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14144 7228 14184 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14144 7140 14184 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14144 7052 14184 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14144 6964 14184 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14063 10111 14103 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14063 10027 14103 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14063 9943 14103 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14063 7580 14103 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14063 7492 14103 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14063 7404 14103 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14063 7316 14103 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14063 7228 14103 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14063 7140 14103 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14063 7052 14103 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 14063 6964 14103 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13982 10111 14022 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13982 10027 14022 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13982 9943 14022 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13982 7580 14022 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13982 7492 14022 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13982 7404 14022 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13982 7316 14022 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13982 7228 14022 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13982 7140 14022 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13982 7052 14022 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13982 6964 14022 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13901 10111 13941 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13901 10027 13941 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13901 9943 13941 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13901 7580 13941 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13901 7492 13941 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13901 7404 13941 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13901 7316 13941 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13901 7228 13941 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13901 7140 13941 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13901 7052 13941 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13901 6964 13941 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13820 10111 13860 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13820 10027 13860 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13820 9943 13860 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13820 7580 13860 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13820 7492 13860 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13820 7404 13860 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13820 7316 13860 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13820 7228 13860 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13820 7140 13860 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13820 7052 13860 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13820 6964 13860 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13739 10111 13779 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13739 10027 13779 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13739 9943 13779 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13739 7580 13779 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13739 7492 13779 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13739 7404 13779 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13739 7316 13779 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13739 7228 13779 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13739 7140 13779 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13739 7052 13779 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13739 6964 13779 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13658 10111 13698 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13658 10027 13698 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13658 9943 13698 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13658 7580 13698 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13658 7492 13698 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13658 7404 13698 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13658 7316 13698 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13658 7228 13698 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13658 7140 13698 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13658 7052 13698 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13658 6964 13698 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13577 10111 13617 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13577 10027 13617 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13577 9943 13617 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13577 7580 13617 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13577 7492 13617 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13577 7404 13617 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13577 7316 13617 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13577 7228 13617 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13577 7140 13617 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13577 7052 13617 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13577 6964 13617 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13496 10111 13536 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13496 10027 13536 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13496 9943 13536 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13496 7580 13536 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13496 7492 13536 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13496 7404 13536 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13496 7316 13536 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13496 7228 13536 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13496 7140 13536 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13496 7052 13536 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13496 6964 13536 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13415 10111 13455 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13415 10027 13455 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13415 9943 13455 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13415 7580 13455 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13415 7492 13455 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13415 7404 13455 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13415 7316 13455 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13415 7228 13455 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13415 7140 13455 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13415 7052 13455 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13415 6964 13455 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13334 10111 13374 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13334 10027 13374 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13334 9943 13374 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13334 7580 13374 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13334 7492 13374 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13334 7404 13374 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13334 7316 13374 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13334 7228 13374 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13334 7140 13374 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13334 7052 13374 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13334 6964 13374 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13253 10111 13293 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13253 10027 13293 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13253 9943 13293 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13253 7580 13293 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13253 7492 13293 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13253 7404 13293 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13253 7316 13293 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13253 7228 13293 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13253 7140 13293 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13253 7052 13293 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13253 6964 13293 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13172 10111 13212 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13172 10027 13212 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13172 9943 13212 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13172 7580 13212 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13172 7492 13212 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13172 7404 13212 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13172 7316 13212 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13172 7228 13212 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13172 7140 13212 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13172 7052 13212 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13172 6964 13212 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13091 10111 13131 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13091 10027 13131 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13091 9943 13131 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13091 7580 13131 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13091 7492 13131 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13091 7404 13131 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13091 7316 13131 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13091 7228 13131 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13091 7140 13131 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13091 7052 13131 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13091 6964 13131 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13010 10111 13050 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13010 10027 13050 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13010 9943 13050 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13010 7580 13050 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13010 7492 13050 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13010 7404 13050 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13010 7316 13050 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13010 7228 13050 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13010 7140 13050 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13010 7052 13050 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 13010 6964 13050 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12929 10111 12969 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12929 10027 12969 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12929 9943 12969 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12929 7580 12969 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12929 7492 12969 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12929 7404 12969 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12929 7316 12969 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12929 7228 12969 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12929 7140 12969 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12929 7052 12969 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12929 6964 12969 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12848 10111 12888 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12848 10027 12888 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12848 9943 12888 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12848 7580 12888 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12848 7492 12888 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12848 7404 12888 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12848 7316 12888 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12848 7228 12888 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12848 7140 12888 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12848 7052 12888 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12848 6964 12888 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12767 10111 12807 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12767 10027 12807 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12767 9943 12807 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12767 7580 12807 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12767 7492 12807 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12767 7404 12807 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12767 7316 12807 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12767 7228 12807 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12767 7140 12807 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12767 7052 12807 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12767 6964 12807 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12686 10111 12726 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12686 10027 12726 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12686 9943 12726 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12686 7580 12726 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12686 7492 12726 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12686 7404 12726 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12686 7316 12726 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12686 7228 12726 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12686 7140 12726 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12686 7052 12726 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12686 6964 12726 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12605 10111 12645 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12605 10027 12645 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12605 9943 12645 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12605 7580 12645 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12605 7492 12645 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12605 7404 12645 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12605 7316 12645 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12605 7228 12645 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12605 7140 12645 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12605 7052 12645 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12605 6964 12645 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12524 10111 12564 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12524 10027 12564 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12524 9943 12564 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12524 7580 12564 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12524 7492 12564 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12524 7404 12564 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12524 7316 12564 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12524 7228 12564 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12524 7140 12564 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12524 7052 12564 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12524 6964 12564 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12443 10111 12483 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12443 10027 12483 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12443 9943 12483 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12443 7580 12483 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12443 7492 12483 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12443 7404 12483 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12443 7316 12483 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12443 7228 12483 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12443 7140 12483 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12443 7052 12483 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12443 6964 12483 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12362 10111 12402 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12362 10027 12402 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12362 9943 12402 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12362 7580 12402 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12362 7492 12402 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12362 7404 12402 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12362 7316 12402 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12362 7228 12402 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12362 7140 12402 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12362 7052 12402 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12362 6964 12402 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12281 10111 12321 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12281 10027 12321 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12281 9943 12321 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12281 7580 12321 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12281 7492 12321 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12281 7404 12321 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12281 7316 12321 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12281 7228 12321 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12281 7140 12321 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12281 7052 12321 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12281 6964 12321 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12200 10111 12240 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12200 10027 12240 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12200 9943 12240 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12200 7580 12240 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12200 7492 12240 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12200 7404 12240 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12200 7316 12240 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12200 7228 12240 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12200 7140 12240 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12200 7052 12240 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12200 6964 12240 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12119 10111 12159 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12119 10027 12159 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12119 9943 12159 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12119 7580 12159 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12119 7492 12159 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12119 7404 12159 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12119 7316 12159 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12119 7228 12159 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12119 7140 12159 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12119 7052 12159 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12119 6964 12159 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12038 10111 12078 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12038 10027 12078 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12038 9943 12078 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12038 7580 12078 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12038 7492 12078 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12038 7404 12078 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12038 7316 12078 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12038 7228 12078 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12038 7140 12078 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12038 7052 12078 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 12038 6964 12078 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11957 10111 11997 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11957 10027 11997 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11957 9943 11997 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11957 7580 11997 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11957 7492 11997 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11957 7404 11997 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11957 7316 11997 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11957 7228 11997 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11957 7140 11997 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11957 7052 11997 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11957 6964 11997 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11876 10111 11916 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11876 10027 11916 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11876 9943 11916 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11876 7580 11916 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11876 7492 11916 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11876 7404 11916 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11876 7316 11916 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11876 7228 11916 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11876 7140 11916 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11876 7052 11916 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11876 6964 11916 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11795 10111 11835 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11795 10027 11835 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11795 9943 11835 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11795 7580 11835 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11795 7492 11835 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11795 7404 11835 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11795 7316 11835 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11795 7228 11835 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11795 7140 11835 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11795 7052 11835 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11795 6964 11835 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11714 10111 11754 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11714 10027 11754 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11714 9943 11754 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11714 7580 11754 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11714 7492 11754 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11714 7404 11754 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11714 7316 11754 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11714 7228 11754 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11714 7140 11754 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11714 7052 11754 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11714 6964 11754 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11633 10111 11673 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11633 10027 11673 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11633 9943 11673 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11633 7580 11673 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11633 7492 11673 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11633 7404 11673 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11633 7316 11673 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11633 7228 11673 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11633 7140 11673 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11633 7052 11673 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11633 6964 11673 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11552 10111 11592 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11552 10027 11592 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11552 9943 11592 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11552 7580 11592 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11552 7492 11592 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11552 7404 11592 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11552 7316 11592 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11552 7228 11592 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11552 7140 11592 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11552 7052 11592 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11552 6964 11592 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11471 10111 11511 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11471 10027 11511 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11471 9943 11511 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11471 7580 11511 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11471 7492 11511 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11471 7404 11511 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11471 7316 11511 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11471 7228 11511 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11471 7140 11511 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11471 7052 11511 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11471 6964 11511 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11390 10111 11430 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11390 10027 11430 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11390 9943 11430 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11390 7580 11430 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11390 7492 11430 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11390 7404 11430 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11390 7316 11430 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11390 7228 11430 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11390 7140 11430 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11390 7052 11430 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11390 6964 11430 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11309 10111 11349 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11309 10027 11349 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11309 9943 11349 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11309 7580 11349 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11309 7492 11349 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11309 7404 11349 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11309 7316 11349 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11309 7228 11349 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11309 7140 11349 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11309 7052 11349 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11309 6964 11349 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11228 10111 11268 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11228 10027 11268 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11228 9943 11268 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11228 7580 11268 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11228 7492 11268 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11228 7404 11268 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11228 7316 11268 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11228 7228 11268 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11228 7140 11268 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11228 7052 11268 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11228 6964 11268 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11147 10111 11187 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11147 10027 11187 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11147 9943 11187 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11147 7580 11187 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11147 7492 11187 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11147 7404 11187 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11147 7316 11187 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11147 7228 11187 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11147 7140 11187 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11147 7052 11187 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11147 6964 11187 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11066 10111 11106 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11066 10027 11106 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11066 9943 11106 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11066 7580 11106 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11066 7492 11106 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11066 7404 11106 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11066 7316 11106 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11066 7228 11106 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11066 7140 11106 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11066 7052 11106 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 11066 6964 11106 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10985 10111 11025 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10985 10027 11025 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10985 9943 11025 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10985 7580 11025 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10985 7492 11025 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10985 7404 11025 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10985 7316 11025 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10985 7228 11025 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10985 7140 11025 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10985 7052 11025 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10985 6964 11025 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10904 10111 10944 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10904 10027 10944 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10904 9943 10944 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10904 7580 10944 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10904 7492 10944 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10904 7404 10944 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10904 7316 10944 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10904 7228 10944 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10904 7140 10944 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10904 7052 10944 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10904 6964 10944 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10823 10111 10863 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10823 10027 10863 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10823 9943 10863 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10823 7580 10863 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10823 7492 10863 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10823 7404 10863 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10823 7316 10863 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10823 7228 10863 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10823 7140 10863 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10823 7052 10863 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10823 6964 10863 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10742 10111 10782 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10742 10027 10782 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10742 9943 10782 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10742 7580 10782 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10742 7492 10782 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10742 7404 10782 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10742 7316 10782 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10742 7228 10782 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10742 7140 10782 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10742 7052 10782 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10742 6964 10782 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10661 10111 10701 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10661 10027 10701 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10661 9943 10701 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10661 7580 10701 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10661 7492 10701 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10661 7404 10701 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10661 7316 10701 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10661 7228 10701 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10661 7140 10701 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10661 7052 10701 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10661 6964 10701 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10579 10111 10619 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10579 10027 10619 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10579 9943 10619 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10579 7580 10619 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10579 7492 10619 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10579 7404 10619 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10579 7316 10619 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10579 7228 10619 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10579 7140 10619 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10579 7052 10619 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10579 6964 10619 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10497 10111 10537 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10497 10027 10537 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10497 9943 10537 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10497 7580 10537 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10497 7492 10537 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10497 7404 10537 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10497 7316 10537 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10497 7228 10537 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10497 7140 10537 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10497 7052 10537 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10497 6964 10537 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10415 10111 10455 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10415 10027 10455 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10415 9943 10455 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10415 7580 10455 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10415 7492 10455 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10415 7404 10455 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10415 7316 10455 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10415 7228 10455 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10415 7140 10455 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10415 7052 10455 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10415 6964 10455 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10333 10111 10373 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10333 10027 10373 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10333 9943 10373 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10333 7580 10373 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10333 7492 10373 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10333 7404 10373 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10333 7316 10373 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10333 7228 10373 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10333 7140 10373 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10333 7052 10373 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10333 6964 10373 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10251 10111 10291 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10251 10027 10291 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10251 9943 10291 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10251 7580 10291 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10251 7492 10291 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10251 7404 10291 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10251 7316 10291 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10251 7228 10291 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10251 7140 10291 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10251 7052 10291 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10251 6964 10291 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10169 10111 10209 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10169 10027 10209 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10169 9943 10209 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10169 7580 10209 7620 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10169 7492 10209 7532 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10169 7404 10209 7444 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10169 7316 10209 7356 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10169 7228 10209 7268 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10169 7140 10209 7180 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10169 7052 10209 7092 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10169 6964 10209 7004 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4822 10111 4862 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4822 10027 4862 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4822 9943 4862 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4810 7568 4874 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4810 7568 4874 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4810 7480 4874 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4810 7480 4874 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4810 7392 4874 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4810 7392 4874 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4810 7304 4874 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4810 7304 4874 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4810 7216 4874 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4810 7216 4874 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4810 7128 4874 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4810 7128 4874 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4810 7040 4874 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4810 7040 4874 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4810 6952 4874 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4810 6952 4874 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4741 10111 4781 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4741 10027 4781 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4741 9943 4781 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4729 7568 4793 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4729 7568 4793 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4729 7480 4793 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4729 7480 4793 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4729 7392 4793 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4729 7392 4793 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4729 7304 4793 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4729 7304 4793 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4729 7216 4793 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4729 7216 4793 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4729 7128 4793 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4729 7128 4793 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4729 7040 4793 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4729 7040 4793 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4729 6952 4793 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4729 6952 4793 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4660 10111 4700 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4660 10027 4700 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4660 9943 4700 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4648 7568 4712 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4648 7568 4712 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4648 7480 4712 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4648 7480 4712 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4648 7392 4712 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4648 7392 4712 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4648 7304 4712 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4648 7304 4712 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4648 7216 4712 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4648 7216 4712 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4648 7128 4712 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4648 7128 4712 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4648 7040 4712 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4648 7040 4712 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4648 6952 4712 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4648 6952 4712 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4579 10111 4619 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4579 10027 4619 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4579 9943 4619 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4567 7568 4631 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4567 7568 4631 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4567 7480 4631 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4567 7480 4631 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4567 7392 4631 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4567 7392 4631 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4567 7304 4631 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4567 7304 4631 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4567 7216 4631 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4567 7216 4631 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4567 7128 4631 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4567 7128 4631 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4567 7040 4631 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4567 7040 4631 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4567 6952 4631 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4567 6952 4631 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4498 10111 4538 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4498 10027 4538 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4498 9943 4538 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4486 7568 4550 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4486 7568 4550 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4486 7480 4550 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4486 7480 4550 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4486 7392 4550 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4486 7392 4550 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4486 7304 4550 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4486 7304 4550 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4486 7216 4550 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4486 7216 4550 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4486 7128 4550 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4486 7128 4550 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4486 7040 4550 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4486 7040 4550 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4486 6952 4550 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4486 6952 4550 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4417 10111 4457 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4417 10027 4457 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4417 9943 4457 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4405 7568 4469 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4405 7568 4469 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4405 7480 4469 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4405 7480 4469 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4405 7392 4469 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4405 7392 4469 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4405 7304 4469 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4405 7304 4469 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4405 7216 4469 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4405 7216 4469 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4405 7128 4469 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4405 7128 4469 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4405 7040 4469 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4405 7040 4469 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4405 6952 4469 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4405 6952 4469 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4336 10111 4376 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4336 10027 4376 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4336 9943 4376 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4324 7568 4388 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4324 7568 4388 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4324 7480 4388 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4324 7480 4388 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4324 7392 4388 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4324 7392 4388 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4324 7304 4388 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4324 7304 4388 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4324 7216 4388 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4324 7216 4388 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4324 7128 4388 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4324 7128 4388 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4324 7040 4388 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4324 7040 4388 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4324 6952 4388 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4324 6952 4388 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4255 10111 4295 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4255 10027 4295 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4255 9943 4295 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4243 7568 4307 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4243 7568 4307 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4243 7480 4307 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4243 7480 4307 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4243 7392 4307 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4243 7392 4307 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4243 7304 4307 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4243 7304 4307 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4243 7216 4307 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4243 7216 4307 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4243 7128 4307 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4243 7128 4307 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4243 7040 4307 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4243 7040 4307 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4243 6952 4307 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4243 6952 4307 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4174 10111 4214 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4174 10027 4214 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4174 9943 4214 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4162 7568 4226 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4162 7568 4226 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4162 7480 4226 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4162 7480 4226 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4162 7392 4226 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4162 7392 4226 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4162 7304 4226 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4162 7304 4226 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4162 7216 4226 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4162 7216 4226 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4162 7128 4226 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4162 7128 4226 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4162 7040 4226 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4162 7040 4226 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4162 6952 4226 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4162 6952 4226 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4093 10111 4133 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4093 10027 4133 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4093 9943 4133 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4081 7568 4145 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4081 7568 4145 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4081 7480 4145 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4081 7480 4145 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4081 7392 4145 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4081 7392 4145 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4081 7304 4145 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4081 7304 4145 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4081 7216 4145 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4081 7216 4145 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4081 7128 4145 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4081 7128 4145 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4081 7040 4145 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4081 7040 4145 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4081 6952 4145 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4081 6952 4145 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4012 10111 4052 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4012 10027 4052 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4012 9943 4052 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4000 7568 4064 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4000 7568 4064 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4000 7480 4064 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4000 7480 4064 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4000 7392 4064 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4000 7392 4064 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4000 7304 4064 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4000 7304 4064 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4000 7216 4064 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4000 7216 4064 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4000 7128 4064 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4000 7128 4064 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4000 7040 4064 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4000 7040 4064 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 4000 6952 4064 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 4000 6952 4064 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3931 10111 3971 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3931 10027 3971 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3931 9943 3971 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3919 7568 3983 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3919 7568 3983 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3919 7480 3983 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3919 7480 3983 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3919 7392 3983 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3919 7392 3983 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3919 7304 3983 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3919 7304 3983 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3919 7216 3983 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3919 7216 3983 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3919 7128 3983 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3919 7128 3983 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3919 7040 3983 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3919 7040 3983 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3919 6952 3983 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3919 6952 3983 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3850 10111 3890 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3850 10027 3890 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3850 9943 3890 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3838 7568 3902 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3838 7568 3902 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3838 7480 3902 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3838 7480 3902 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3838 7392 3902 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3838 7392 3902 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3838 7304 3902 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3838 7304 3902 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3838 7216 3902 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3838 7216 3902 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3838 7128 3902 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3838 7128 3902 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3838 7040 3902 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3838 7040 3902 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3838 6952 3902 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3838 6952 3902 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3769 10111 3809 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3769 10027 3809 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3769 9943 3809 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3757 7568 3821 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3757 7568 3821 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3757 7480 3821 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3757 7480 3821 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3757 7392 3821 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3757 7392 3821 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3757 7304 3821 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3757 7304 3821 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3757 7216 3821 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3757 7216 3821 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3757 7128 3821 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3757 7128 3821 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3757 7040 3821 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3757 7040 3821 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3757 6952 3821 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3757 6952 3821 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3688 10111 3728 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3688 10027 3728 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3688 9943 3728 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3676 7568 3740 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3676 7568 3740 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3676 7480 3740 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3676 7480 3740 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3676 7392 3740 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3676 7392 3740 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3676 7304 3740 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3676 7304 3740 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3676 7216 3740 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3676 7216 3740 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3676 7128 3740 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3676 7128 3740 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3676 7040 3740 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3676 7040 3740 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3676 6952 3740 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3676 6952 3740 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3607 10111 3647 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3607 10027 3647 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3607 9943 3647 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3595 7568 3659 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3595 7568 3659 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3595 7480 3659 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3595 7480 3659 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3595 7392 3659 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3595 7392 3659 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3595 7304 3659 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3595 7304 3659 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3595 7216 3659 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3595 7216 3659 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3595 7128 3659 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3595 7128 3659 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3595 7040 3659 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3595 7040 3659 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3595 6952 3659 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3595 6952 3659 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3526 10111 3566 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3526 10027 3566 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3526 9943 3566 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3514 7568 3578 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3514 7568 3578 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3514 7480 3578 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3514 7480 3578 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3514 7392 3578 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3514 7392 3578 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3514 7304 3578 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3514 7304 3578 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3514 7216 3578 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3514 7216 3578 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3514 7128 3578 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3514 7128 3578 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3514 7040 3578 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3514 7040 3578 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3514 6952 3578 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3514 6952 3578 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3445 10111 3485 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3445 10027 3485 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3445 9943 3485 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3433 7568 3497 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3433 7568 3497 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3433 7480 3497 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3433 7480 3497 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3433 7392 3497 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3433 7392 3497 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3433 7304 3497 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3433 7304 3497 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3433 7216 3497 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3433 7216 3497 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3433 7128 3497 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3433 7128 3497 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3433 7040 3497 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3433 7040 3497 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3433 6952 3497 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3433 6952 3497 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3364 10111 3404 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3364 10027 3404 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3364 9943 3404 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3352 7568 3416 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3352 7568 3416 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3352 7480 3416 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3352 7480 3416 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3352 7392 3416 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3352 7392 3416 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3352 7304 3416 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3352 7304 3416 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3352 7216 3416 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3352 7216 3416 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3352 7128 3416 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3352 7128 3416 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3352 7040 3416 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3352 7040 3416 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3352 6952 3416 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3352 6952 3416 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3283 10111 3323 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3283 10027 3323 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3283 9943 3323 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3271 7568 3335 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3271 7568 3335 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3271 7480 3335 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3271 7480 3335 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3271 7392 3335 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3271 7392 3335 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3271 7304 3335 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3271 7304 3335 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3271 7216 3335 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3271 7216 3335 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3271 7128 3335 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3271 7128 3335 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3271 7040 3335 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3271 7040 3335 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3271 6952 3335 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3271 6952 3335 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3202 10111 3242 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3202 10027 3242 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3202 9943 3242 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3190 7568 3254 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3190 7568 3254 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3190 7480 3254 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3190 7480 3254 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3190 7392 3254 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3190 7392 3254 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3190 7304 3254 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3190 7304 3254 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3190 7216 3254 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3190 7216 3254 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3190 7128 3254 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3190 7128 3254 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3190 7040 3254 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3190 7040 3254 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3190 6952 3254 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3190 6952 3254 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3121 10111 3161 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3121 10027 3161 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3121 9943 3161 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3109 7568 3173 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3109 7568 3173 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3109 7480 3173 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3109 7480 3173 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3109 7392 3173 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3109 7392 3173 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3109 7304 3173 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3109 7304 3173 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3109 7216 3173 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3109 7216 3173 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3109 7128 3173 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3109 7128 3173 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3109 7040 3173 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3109 7040 3173 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3109 6952 3173 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3109 6952 3173 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3040 10111 3080 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3040 10027 3080 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3040 9943 3080 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3028 7568 3092 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3028 7568 3092 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3028 7480 3092 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3028 7480 3092 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3028 7392 3092 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3028 7392 3092 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3028 7304 3092 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3028 7304 3092 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3028 7216 3092 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3028 7216 3092 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3028 7128 3092 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3028 7128 3092 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3028 7040 3092 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3028 7040 3092 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 3028 6952 3092 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 3028 6952 3092 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2959 10111 2999 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2959 10027 2999 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2959 9943 2999 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2947 7568 3011 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2947 7568 3011 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2947 7480 3011 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2947 7480 3011 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2947 7392 3011 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2947 7392 3011 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2947 7304 3011 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2947 7304 3011 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2947 7216 3011 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2947 7216 3011 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2947 7128 3011 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2947 7128 3011 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2947 7040 3011 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2947 7040 3011 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2947 6952 3011 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2947 6952 3011 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2878 10111 2918 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2878 10027 2918 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2878 9943 2918 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2866 7568 2930 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2866 7568 2930 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2866 7480 2930 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2866 7480 2930 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2866 7392 2930 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2866 7392 2930 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2866 7304 2930 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2866 7304 2930 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2866 7216 2930 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2866 7216 2930 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2866 7128 2930 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2866 7128 2930 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2866 7040 2930 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2866 7040 2930 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2866 6952 2930 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2866 6952 2930 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2797 10111 2837 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2797 10027 2837 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2797 9943 2837 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2785 7568 2849 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2785 7568 2849 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2785 7480 2849 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2785 7480 2849 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2785 7392 2849 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2785 7392 2849 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2785 7304 2849 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2785 7304 2849 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2785 7216 2849 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2785 7216 2849 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2785 7128 2849 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2785 7128 2849 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2785 7040 2849 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2785 7040 2849 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2785 6952 2849 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2785 6952 2849 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2716 10111 2756 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2716 10027 2756 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2716 9943 2756 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2704 7568 2768 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2704 7568 2768 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2704 7480 2768 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2704 7480 2768 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2704 7392 2768 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2704 7392 2768 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2704 7304 2768 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2704 7304 2768 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2704 7216 2768 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2704 7216 2768 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2704 7128 2768 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2704 7128 2768 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2704 7040 2768 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2704 7040 2768 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2704 6952 2768 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2704 6952 2768 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2635 10111 2675 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2635 10027 2675 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2635 9943 2675 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2623 7568 2687 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2623 7568 2687 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2623 7480 2687 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2623 7480 2687 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2623 7392 2687 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2623 7392 2687 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2623 7304 2687 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2623 7304 2687 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2623 7216 2687 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2623 7216 2687 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2623 7128 2687 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2623 7128 2687 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2623 7040 2687 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2623 7040 2687 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2623 6952 2687 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2623 6952 2687 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2554 10111 2594 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2554 10027 2594 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2554 9943 2594 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2542 7568 2606 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2542 7568 2606 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2542 7480 2606 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2542 7480 2606 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2542 7392 2606 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2542 7392 2606 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2542 7304 2606 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2542 7304 2606 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2542 7216 2606 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2542 7216 2606 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2542 7128 2606 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2542 7128 2606 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2542 7040 2606 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2542 7040 2606 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2542 6952 2606 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2542 6952 2606 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2473 10111 2513 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2473 10027 2513 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2473 9943 2513 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2461 7568 2525 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2461 7568 2525 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2461 7480 2525 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2461 7480 2525 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2461 7392 2525 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2461 7392 2525 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2461 7304 2525 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2461 7304 2525 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2461 7216 2525 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2461 7216 2525 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2461 7128 2525 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2461 7128 2525 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2461 7040 2525 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2461 7040 2525 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2461 6952 2525 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2461 6952 2525 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2392 10111 2432 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2392 10027 2432 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2392 9943 2432 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2380 7568 2444 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2380 7568 2444 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2380 7480 2444 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2380 7480 2444 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2380 7392 2444 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2380 7392 2444 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2380 7304 2444 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2380 7304 2444 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2380 7216 2444 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2380 7216 2444 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2380 7128 2444 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2380 7128 2444 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2380 7040 2444 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2380 7040 2444 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2380 6952 2444 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2380 6952 2444 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2311 10111 2351 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2311 10027 2351 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2311 9943 2351 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2299 7568 2363 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2299 7568 2363 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2299 7480 2363 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2299 7480 2363 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2299 7392 2363 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2299 7392 2363 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2299 7304 2363 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2299 7304 2363 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2299 7216 2363 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2299 7216 2363 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2299 7128 2363 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2299 7128 2363 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2299 7040 2363 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2299 7040 2363 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2299 6952 2363 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2299 6952 2363 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2230 10111 2270 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2230 10027 2270 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2230 9943 2270 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2218 7568 2282 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2218 7568 2282 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2218 7480 2282 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2218 7480 2282 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2218 7392 2282 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2218 7392 2282 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2218 7304 2282 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2218 7304 2282 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2218 7216 2282 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2218 7216 2282 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2218 7128 2282 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2218 7128 2282 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2218 7040 2282 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2218 7040 2282 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2218 6952 2282 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2218 6952 2282 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2149 10111 2189 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2149 10027 2189 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2149 9943 2189 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2137 7568 2201 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2137 7568 2201 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2137 7480 2201 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2137 7480 2201 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2137 7392 2201 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2137 7392 2201 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2137 7304 2201 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2137 7304 2201 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2137 7216 2201 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2137 7216 2201 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2137 7128 2201 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2137 7128 2201 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2137 7040 2201 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2137 7040 2201 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2137 6952 2201 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2137 6952 2201 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2068 10111 2108 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2068 10027 2108 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2068 9943 2108 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2056 7568 2120 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2056 7568 2120 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2056 7480 2120 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2056 7480 2120 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2056 7392 2120 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2056 7392 2120 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2056 7304 2120 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2056 7304 2120 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2056 7216 2120 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2056 7216 2120 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2056 7128 2120 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2056 7128 2120 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2056 7040 2120 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2056 7040 2120 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 2056 6952 2120 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 2056 6952 2120 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1987 10111 2027 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1987 10027 2027 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1987 9943 2027 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1975 7568 2039 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1975 7568 2039 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1975 7480 2039 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1975 7480 2039 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1975 7392 2039 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1975 7392 2039 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1975 7304 2039 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1975 7304 2039 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1975 7216 2039 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1975 7216 2039 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1975 7128 2039 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1975 7128 2039 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1975 7040 2039 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1975 7040 2039 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1975 6952 2039 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1975 6952 2039 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1906 10111 1946 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1906 10027 1946 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1906 9943 1946 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1894 7568 1958 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1894 7568 1958 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1894 7480 1958 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1894 7480 1958 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1894 7392 1958 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1894 7392 1958 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1894 7304 1958 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1894 7304 1958 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1894 7216 1958 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1894 7216 1958 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1894 7128 1958 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1894 7128 1958 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1894 7040 1958 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1894 7040 1958 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1894 6952 1958 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1894 6952 1958 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1825 10111 1865 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1825 10027 1865 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1825 9943 1865 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1813 7568 1877 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1813 7568 1877 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1813 7480 1877 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1813 7480 1877 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1813 7392 1877 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1813 7392 1877 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1813 7304 1877 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1813 7304 1877 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1813 7216 1877 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1813 7216 1877 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1813 7128 1877 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1813 7128 1877 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1813 7040 1877 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1813 7040 1877 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1813 6952 1877 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1813 6952 1877 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1744 10111 1784 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1744 10027 1784 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1744 9943 1784 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1732 7568 1796 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1732 7568 1796 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1732 7480 1796 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1732 7480 1796 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1732 7392 1796 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1732 7392 1796 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1732 7304 1796 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1732 7304 1796 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1732 7216 1796 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1732 7216 1796 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1732 7128 1796 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1732 7128 1796 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1732 7040 1796 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1732 7040 1796 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1732 6952 1796 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1732 6952 1796 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1663 10111 1703 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1663 10027 1703 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1663 9943 1703 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1651 7568 1715 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1651 7568 1715 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1651 7480 1715 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1651 7480 1715 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1651 7392 1715 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1651 7392 1715 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1651 7304 1715 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1651 7304 1715 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1651 7216 1715 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1651 7216 1715 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1651 7128 1715 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1651 7128 1715 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1651 7040 1715 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1651 7040 1715 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1651 6952 1715 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1651 6952 1715 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1582 10111 1622 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1582 10027 1622 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1582 9943 1622 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1570 7568 1634 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1570 7568 1634 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1570 7480 1634 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1570 7480 1634 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1570 7392 1634 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1570 7392 1634 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1570 7304 1634 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1570 7304 1634 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1570 7216 1634 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1570 7216 1634 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1570 7128 1634 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1570 7128 1634 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1570 7040 1634 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1570 7040 1634 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1570 6952 1634 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1570 6952 1634 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1501 10111 1541 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1501 10027 1541 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1501 9943 1541 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1489 7568 1553 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1489 7568 1553 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1489 7480 1553 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1489 7480 1553 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1489 7392 1553 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1489 7392 1553 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1489 7304 1553 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1489 7304 1553 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1489 7216 1553 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1489 7216 1553 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1489 7128 1553 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1489 7128 1553 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1489 7040 1553 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1489 7040 1553 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1489 6952 1553 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1489 6952 1553 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1420 10111 1460 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1420 10027 1460 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1420 9943 1460 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1408 7568 1472 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1408 7568 1472 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1408 7480 1472 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1408 7480 1472 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1408 7392 1472 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1408 7392 1472 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1408 7304 1472 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1408 7304 1472 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1408 7216 1472 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1408 7216 1472 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1408 7128 1472 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1408 7128 1472 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1408 7040 1472 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1408 7040 1472 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1408 6952 1472 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1408 6952 1472 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1339 10111 1379 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1339 10027 1379 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1339 9943 1379 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1327 7568 1391 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1327 7568 1391 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1327 7480 1391 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1327 7480 1391 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1327 7392 1391 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1327 7392 1391 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1327 7304 1391 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1327 7304 1391 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1327 7216 1391 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1327 7216 1391 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1327 7128 1391 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1327 7128 1391 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1327 7040 1391 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1327 7040 1391 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1327 6952 1391 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1327 6952 1391 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1258 10111 1298 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1258 10027 1298 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1258 9943 1298 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1246 7568 1310 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1246 7568 1310 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1246 7480 1310 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1246 7480 1310 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1246 7392 1310 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1246 7392 1310 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1246 7304 1310 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1246 7304 1310 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1246 7216 1310 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1246 7216 1310 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1246 7128 1310 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1246 7128 1310 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1246 7040 1310 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1246 7040 1310 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1246 6952 1310 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1246 6952 1310 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1177 10111 1217 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1177 10027 1217 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1177 9943 1217 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1165 7568 1229 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1165 7568 1229 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1165 7480 1229 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1165 7480 1229 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1165 7392 1229 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1165 7392 1229 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1165 7304 1229 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1165 7304 1229 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1165 7216 1229 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1165 7216 1229 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1165 7128 1229 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1165 7128 1229 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1165 7040 1229 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1165 7040 1229 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1165 6952 1229 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1165 6952 1229 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1096 10111 1136 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1096 10027 1136 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1096 9943 1136 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1084 7568 1148 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1084 7568 1148 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1084 7480 1148 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1084 7480 1148 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1084 7392 1148 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1084 7392 1148 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1084 7304 1148 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1084 7304 1148 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1084 7216 1148 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1084 7216 1148 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1084 7128 1148 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1084 7128 1148 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1084 7040 1148 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1084 7040 1148 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1084 6952 1148 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1084 6952 1148 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1015 10111 1055 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1015 10027 1055 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1015 9943 1055 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1003 7568 1067 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1003 7568 1067 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1003 7480 1067 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1003 7480 1067 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1003 7392 1067 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1003 7392 1067 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1003 7304 1067 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1003 7304 1067 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1003 7216 1067 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1003 7216 1067 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1003 7128 1067 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1003 7128 1067 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1003 7040 1067 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1003 7040 1067 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 1003 6952 1067 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 1003 6952 1067 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 934 10111 974 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 934 10027 974 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 934 9943 974 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 922 7568 986 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 922 7568 986 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 922 7480 986 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 922 7480 986 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 922 7392 986 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 922 7392 986 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 922 7304 986 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 922 7304 986 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 922 7216 986 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 922 7216 986 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 922 7128 986 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 922 7128 986 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 922 7040 986 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 922 7040 986 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 922 6952 986 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 922 6952 986 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 853 10111 893 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 853 10027 893 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 853 9943 893 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 841 7568 905 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 841 7568 905 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 841 7480 905 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 841 7480 905 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 841 7392 905 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 841 7392 905 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 841 7304 905 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 841 7304 905 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 841 7216 905 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 841 7216 905 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 841 7128 905 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 841 7128 905 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 841 7040 905 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 841 7040 905 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 841 6952 905 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 841 6952 905 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 772 10111 812 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 772 10027 812 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 772 9943 812 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 760 7568 824 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 760 7568 824 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 760 7480 824 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 760 7480 824 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 760 7392 824 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 760 7392 824 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 760 7304 824 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 760 7304 824 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 760 7216 824 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 760 7216 824 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 760 7128 824 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 760 7128 824 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 760 7040 824 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 760 7040 824 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 760 6952 824 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 760 6952 824 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 691 10111 731 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 691 10027 731 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 691 9943 731 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 679 7568 743 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 679 7568 743 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 679 7480 743 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 679 7480 743 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 679 7392 743 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 679 7392 743 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 679 7304 743 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 679 7304 743 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 679 7216 743 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 679 7216 743 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 679 7128 743 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 679 7128 743 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 679 7040 743 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 679 7040 743 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 679 6952 743 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 679 6952 743 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 610 10111 650 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 610 10027 650 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 610 9943 650 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 598 7568 662 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 598 7568 662 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 598 7480 662 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 598 7480 662 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 598 7392 662 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 598 7392 662 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 598 7304 662 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 598 7304 662 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 598 7216 662 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 598 7216 662 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 598 7128 662 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 598 7128 662 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 598 7040 662 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 598 7040 662 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 598 6952 662 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 598 6952 662 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 528 10111 568 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 528 10027 568 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 528 9943 568 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 516 7568 580 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 516 7568 580 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 516 7480 580 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 516 7480 580 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 516 7392 580 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 516 7392 580 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 516 7304 580 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 516 7304 580 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 516 7216 580 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 516 7216 580 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 516 7128 580 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 516 7128 580 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 516 7040 580 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 516 7040 580 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 516 6952 580 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 516 6952 580 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 446 10111 486 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 446 10027 486 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 446 9943 486 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 434 7568 498 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 434 7568 498 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 434 7480 498 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 434 7480 498 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 434 7392 498 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 434 7392 498 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 434 7304 498 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 434 7304 498 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 434 7216 498 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 434 7216 498 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 434 7128 498 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 434 7128 498 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 434 7040 498 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 434 7040 498 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 434 6952 498 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 434 6952 498 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 364 10111 404 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 364 10027 404 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 364 9943 404 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 352 7568 416 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 352 7568 416 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 352 7480 416 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 352 7480 416 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 352 7392 416 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 352 7392 416 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 352 7304 416 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 352 7304 416 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 352 7216 416 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 352 7216 416 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 352 7128 416 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 352 7128 416 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 352 7040 416 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 352 7040 416 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 352 6952 416 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 352 6952 416 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 282 10111 322 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 282 10027 322 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 282 9943 322 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 270 7568 334 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 270 7568 334 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 270 7480 334 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 270 7480 334 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 270 7392 334 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 270 7392 334 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 270 7304 334 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 270 7304 334 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 270 7216 334 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 270 7216 334 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 270 7128 334 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 270 7128 334 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 270 7040 334 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 270 7040 334 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 270 6952 334 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 270 6952 334 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 200 10111 240 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 200 10027 240 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 200 9943 240 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 188 7568 252 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 188 7480 252 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 188 7392 252 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 188 7304 252 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 188 7216 252 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 188 7128 252 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 188 7040 252 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 188 6952 252 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 118 10111 158 10151 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 118 10027 158 10067 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 118 9943 158 9983 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 106 7568 170 7632 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 106 7480 170 7544 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 106 7392 170 7456 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 106 7304 170 7368 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 106 7216 170 7280 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 106 7128 170 7192 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 106 7040 170 7104 6 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 106 6952 170 7016 6 VSSA
port 2 nsew ground bidirectional
rlabel metal5 s 0 27 254 1077 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal4 s 0 7 254 1097 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal5 s 14746 7937 15000 8827 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 0 7917 254 8847 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 34757 254 39600 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 4767 254 5697 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 6 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal5 s 0 11267 254 12117 6 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 6 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal4 s 0 11247 254 12137 6 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 VCCD
port 7 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 6 VCCD
port 7 nsew power bidirectional
rlabel metal4 s 0 1377 254 2307 6 VCCD
port 7 nsew power bidirectional
rlabel metal4 s 14746 1377 15000 2307 6 VCCD
port 7 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 0 2587 193 3277 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 6 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 6 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 6 VDDIO
port 9 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 6 VDDIO
port 9 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 6 VDDIO
port 9 nsew power bidirectional
rlabel metal4 s 0 3557 254 4487 6 VDDIO
port 9 nsew power bidirectional
rlabel metal4 s 0 13607 254 18600 6 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 14746 5997 15000 6647 6 VSWITCH
port 10 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 6 VSWITCH
port 10 nsew power bidirectional
rlabel metal4 s 14746 5977 15000 6667 6 VSWITCH
port 10 nsew power bidirectional
rlabel metal4 s 0 5977 254 6667 6 VSWITCH
port 10 nsew power bidirectional
rlabel metal4 s 0 10225 15000 10821 6 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 0 9273 15000 9869 6 AMUXBUS_B
port 12 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 39600
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 25710796
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 25619004
<< end >>
