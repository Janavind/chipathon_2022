magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 834 157 1653 203
rect 1 21 1653 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 435 47 465 131
rect 543 47 573 119
rect 629 47 659 119
rect 724 47 754 131
rect 912 47 942 177
rect 996 47 1026 177
rect 1080 47 1110 177
rect 1175 47 1205 177
rect 1365 47 1395 131
rect 1460 47 1490 177
rect 1545 47 1575 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 435 369 465 497
rect 531 413 561 497
rect 652 413 682 497
rect 724 413 754 497
rect 912 297 942 497
rect 996 297 1026 497
rect 1080 297 1110 497
rect 1175 297 1205 497
rect 1365 369 1395 497
rect 1460 297 1490 497
rect 1545 297 1575 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 119 351 131
rect 299 85 307 119
rect 341 85 351 119
rect 299 47 351 85
rect 381 89 435 131
rect 381 55 391 89
rect 425 55 435 89
rect 381 47 435 55
rect 465 119 515 131
rect 860 133 912 177
rect 674 119 724 131
rect 465 47 543 119
rect 573 107 629 119
rect 573 73 584 107
rect 618 73 629 107
rect 573 47 629 73
rect 659 47 724 119
rect 754 106 806 131
rect 754 72 764 106
rect 798 72 806 106
rect 754 47 806 72
rect 860 99 868 133
rect 902 99 912 133
rect 860 47 912 99
rect 942 47 996 177
rect 1026 89 1080 177
rect 1026 55 1036 89
rect 1070 55 1080 89
rect 1026 47 1080 55
rect 1110 133 1175 177
rect 1110 99 1130 133
rect 1164 99 1175 133
rect 1110 47 1175 99
rect 1205 93 1259 177
rect 1410 131 1460 177
rect 1205 59 1217 93
rect 1251 59 1259 93
rect 1205 47 1259 59
rect 1313 119 1365 131
rect 1313 85 1321 119
rect 1355 85 1365 119
rect 1313 47 1365 85
rect 1395 93 1460 131
rect 1395 59 1416 93
rect 1450 59 1460 93
rect 1395 47 1460 59
rect 1490 129 1545 177
rect 1490 95 1500 129
rect 1534 95 1545 129
rect 1490 47 1545 95
rect 1575 161 1627 177
rect 1575 127 1585 161
rect 1619 127 1627 161
rect 1575 93 1627 127
rect 1575 59 1585 93
rect 1619 59 1627 93
rect 1575 47 1627 59
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 483 351 497
rect 299 449 307 483
rect 341 449 351 483
rect 299 415 351 449
rect 299 381 307 415
rect 341 381 351 415
rect 299 369 351 381
rect 381 485 435 497
rect 381 451 391 485
rect 425 451 435 485
rect 381 417 435 451
rect 381 383 391 417
rect 425 383 435 417
rect 381 369 435 383
rect 465 413 531 497
rect 561 485 652 497
rect 561 451 596 485
rect 630 451 652 485
rect 561 413 652 451
rect 682 413 724 497
rect 754 477 806 497
rect 754 443 764 477
rect 798 443 806 477
rect 754 413 806 443
rect 860 485 912 497
rect 860 451 868 485
rect 902 451 912 485
rect 465 369 515 413
rect 860 297 912 451
rect 942 471 996 497
rect 942 437 952 471
rect 986 437 996 471
rect 942 368 996 437
rect 942 334 952 368
rect 986 334 996 368
rect 942 297 996 334
rect 1026 489 1080 497
rect 1026 455 1036 489
rect 1070 455 1080 489
rect 1026 421 1080 455
rect 1026 387 1036 421
rect 1070 387 1080 421
rect 1026 297 1080 387
rect 1110 477 1175 497
rect 1110 443 1130 477
rect 1164 443 1175 477
rect 1110 409 1175 443
rect 1110 375 1130 409
rect 1164 375 1175 409
rect 1110 297 1175 375
rect 1205 485 1259 497
rect 1205 451 1217 485
rect 1251 451 1259 485
rect 1205 417 1259 451
rect 1205 383 1217 417
rect 1251 383 1259 417
rect 1205 297 1259 383
rect 1313 485 1365 497
rect 1313 451 1321 485
rect 1355 451 1365 485
rect 1313 417 1365 451
rect 1313 383 1321 417
rect 1355 383 1365 417
rect 1313 369 1365 383
rect 1395 485 1460 497
rect 1395 451 1416 485
rect 1450 451 1460 485
rect 1395 417 1460 451
rect 1395 383 1416 417
rect 1450 383 1460 417
rect 1395 369 1460 383
rect 1410 297 1460 369
rect 1490 449 1545 497
rect 1490 415 1500 449
rect 1534 415 1545 449
rect 1490 381 1545 415
rect 1490 347 1500 381
rect 1534 347 1545 381
rect 1490 297 1545 347
rect 1575 485 1627 497
rect 1575 451 1585 485
rect 1619 451 1627 485
rect 1575 417 1627 451
rect 1575 383 1585 417
rect 1619 383 1627 417
rect 1575 349 1627 383
rect 1575 315 1585 349
rect 1619 315 1627 349
rect 1575 297 1627 315
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 85 341 119
rect 391 55 425 89
rect 584 73 618 107
rect 764 72 798 106
rect 868 99 902 133
rect 1036 55 1070 89
rect 1130 99 1164 133
rect 1217 59 1251 93
rect 1321 85 1355 119
rect 1416 59 1450 93
rect 1500 95 1534 129
rect 1585 127 1619 161
rect 1585 59 1619 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 449 341 483
rect 307 381 341 415
rect 391 451 425 485
rect 391 383 425 417
rect 596 451 630 485
rect 764 443 798 477
rect 868 451 902 485
rect 952 437 986 471
rect 952 334 986 368
rect 1036 455 1070 489
rect 1036 387 1070 421
rect 1130 443 1164 477
rect 1130 375 1164 409
rect 1217 451 1251 485
rect 1217 383 1251 417
rect 1321 451 1355 485
rect 1321 383 1355 417
rect 1416 451 1450 485
rect 1416 383 1450 417
rect 1500 415 1534 449
rect 1500 347 1534 381
rect 1585 451 1619 485
rect 1585 383 1619 417
rect 1585 315 1619 349
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 435 497 465 523
rect 531 497 561 523
rect 652 497 682 523
rect 724 497 754 523
rect 912 497 942 523
rect 996 497 1026 523
rect 1080 497 1110 523
rect 1175 497 1205 523
rect 1365 497 1395 523
rect 1460 497 1490 523
rect 1545 497 1575 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 21 264 76 280
rect 163 274 193 363
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 351 241 381 369
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 298 225 381 241
rect 298 191 308 225
rect 342 191 381 225
rect 435 219 465 369
rect 531 337 561 413
rect 652 375 682 413
rect 507 321 561 337
rect 603 365 682 375
rect 603 331 619 365
rect 653 331 682 365
rect 603 321 682 331
rect 724 373 754 413
rect 724 357 812 373
rect 724 323 768 357
rect 802 323 812 357
rect 507 287 517 321
rect 551 287 561 321
rect 507 279 561 287
rect 724 307 812 323
rect 507 271 659 279
rect 531 249 659 271
rect 298 175 381 191
rect 351 131 381 175
rect 424 203 478 219
rect 424 169 434 203
rect 468 169 478 203
rect 424 153 478 169
rect 533 191 587 207
rect 533 157 543 191
rect 577 157 587 191
rect 435 131 465 153
rect 533 141 587 157
rect 543 119 573 141
rect 629 119 659 249
rect 724 131 754 307
rect 1365 354 1395 369
rect 1339 324 1395 354
rect 912 265 942 297
rect 996 265 1026 297
rect 1080 265 1110 297
rect 1175 265 1205 297
rect 1339 265 1369 324
rect 1460 265 1490 297
rect 796 249 942 265
rect 796 215 806 249
rect 840 215 942 249
rect 796 199 942 215
rect 984 249 1038 265
rect 984 215 994 249
rect 1028 215 1038 249
rect 984 199 1038 215
rect 1080 249 1369 265
rect 1080 215 1090 249
rect 1124 215 1369 249
rect 1080 199 1369 215
rect 1431 259 1490 265
rect 1545 259 1575 297
rect 1431 249 1575 259
rect 1431 215 1441 249
rect 1475 215 1575 249
rect 1431 205 1575 215
rect 1431 199 1490 205
rect 912 177 942 199
rect 996 177 1026 199
rect 1080 177 1110 199
rect 1175 177 1205 199
rect 1339 176 1369 199
rect 1460 177 1490 199
rect 1545 177 1575 205
rect 1339 146 1395 176
rect 1365 131 1395 146
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 435 21 465 47
rect 543 21 573 47
rect 629 21 659 47
rect 724 21 754 47
rect 912 21 942 47
rect 996 21 1026 47
rect 1080 21 1110 47
rect 1175 21 1205 47
rect 1365 21 1395 47
rect 1460 21 1490 47
rect 1545 21 1575 47
<< polycont >>
rect 32 230 66 264
rect 134 230 168 264
rect 308 191 342 225
rect 619 331 653 365
rect 768 323 802 357
rect 517 287 551 321
rect 434 169 468 203
rect 543 157 577 191
rect 806 215 840 249
rect 994 215 1028 249
rect 1090 215 1124 249
rect 1441 215 1475 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 17 477 69 493
rect 17 443 35 477
rect 17 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 391 485 454 527
rect 764 485 918 527
rect 1020 489 1070 527
rect 237 443 248 477
rect 17 375 35 409
rect 203 409 248 443
rect 69 375 156 393
rect 17 359 156 375
rect 17 264 66 325
rect 17 230 32 264
rect 17 197 66 230
rect 121 323 156 359
rect 121 289 122 323
rect 121 280 156 289
rect 237 391 248 409
rect 203 357 214 375
rect 203 337 248 357
rect 291 449 307 483
rect 341 449 357 483
rect 291 415 357 449
rect 291 381 307 415
rect 341 381 357 415
rect 121 264 168 280
rect 121 230 134 264
rect 121 214 168 230
rect 121 161 156 214
rect 17 127 156 161
rect 17 119 69 127
rect 17 85 35 119
rect 203 119 237 337
rect 291 333 357 381
rect 425 451 454 485
rect 580 451 596 485
rect 630 451 730 485
rect 391 417 454 451
rect 425 383 454 417
rect 391 367 454 383
rect 494 391 551 401
rect 528 357 551 391
rect 291 299 428 333
rect 292 225 358 265
rect 292 191 308 225
rect 342 191 358 225
rect 394 219 428 299
rect 494 321 551 357
rect 494 287 517 321
rect 494 271 551 287
rect 585 365 653 399
rect 585 331 619 365
rect 585 323 653 331
rect 585 289 586 323
rect 620 289 653 323
rect 585 283 653 289
rect 394 203 468 219
rect 585 207 619 283
rect 696 265 730 451
rect 764 477 868 485
rect 798 451 868 477
rect 902 451 918 485
rect 798 443 918 451
rect 764 427 918 443
rect 952 471 986 487
rect 952 373 986 437
rect 768 368 986 373
rect 1020 455 1036 489
rect 1020 421 1070 455
rect 1020 387 1036 421
rect 1020 371 1070 387
rect 1130 477 1183 493
rect 1164 443 1183 477
rect 1130 409 1183 443
rect 1164 375 1183 409
rect 768 357 952 368
rect 802 334 952 357
rect 802 333 986 334
rect 802 323 1096 333
rect 768 299 1096 323
rect 1130 332 1183 375
rect 1217 485 1271 527
rect 1251 451 1271 485
rect 1217 417 1271 451
rect 1251 383 1271 417
rect 1217 366 1271 383
rect 1305 485 1371 493
rect 1305 451 1321 485
rect 1355 451 1371 485
rect 1305 417 1371 451
rect 1305 383 1321 417
rect 1355 383 1371 417
rect 1130 299 1195 332
rect 1062 265 1096 299
rect 1158 265 1195 299
rect 1305 265 1371 383
rect 1407 485 1466 527
rect 1407 451 1416 485
rect 1450 451 1466 485
rect 1407 417 1466 451
rect 1407 383 1416 417
rect 1450 383 1466 417
rect 1407 367 1466 383
rect 1500 449 1551 493
rect 1534 415 1551 449
rect 1500 381 1551 415
rect 1534 347 1551 381
rect 1500 289 1551 347
rect 1585 485 1639 527
rect 1619 451 1639 485
rect 1585 417 1639 451
rect 1619 383 1639 417
rect 1585 349 1639 383
rect 1619 315 1639 349
rect 1585 299 1639 315
rect 1509 265 1551 289
rect 696 249 840 265
rect 696 233 806 249
rect 394 169 434 203
rect 394 157 468 169
rect 17 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 307 153 468 157
rect 543 191 619 207
rect 577 157 619 191
rect 307 123 428 153
rect 543 141 619 157
rect 666 215 806 233
rect 666 199 840 215
rect 878 249 1028 265
rect 878 215 994 249
rect 878 199 1028 215
rect 1062 249 1124 265
rect 1062 215 1090 249
rect 1062 199 1124 215
rect 307 119 341 123
rect 666 107 700 199
rect 1062 165 1096 199
rect 1158 177 1271 265
rect 1305 249 1475 265
rect 1305 215 1441 249
rect 1305 199 1475 215
rect 1509 211 1639 265
rect 1158 172 1195 177
rect 1148 165 1195 172
rect 307 69 341 85
rect 103 17 169 59
rect 375 55 391 89
rect 425 55 441 89
rect 568 73 584 107
rect 618 73 700 107
rect 748 106 814 165
rect 375 17 441 55
rect 748 72 764 106
rect 798 72 814 106
rect 868 133 1096 165
rect 902 131 1096 133
rect 1130 137 1195 165
rect 1130 133 1190 137
rect 902 99 912 131
rect 868 83 912 99
rect 1164 131 1190 133
rect 1164 99 1182 131
rect 1305 119 1371 199
rect 1509 165 1551 211
rect 1020 89 1096 97
rect 748 17 814 72
rect 1020 55 1036 89
rect 1070 55 1096 89
rect 1130 83 1182 99
rect 1217 93 1271 109
rect 1020 17 1096 55
rect 1251 59 1271 93
rect 1217 17 1271 59
rect 1305 85 1321 119
rect 1355 85 1371 119
rect 1500 129 1551 165
rect 1305 51 1371 85
rect 1405 93 1466 109
rect 1405 59 1416 93
rect 1450 59 1466 93
rect 1405 17 1466 59
rect 1534 95 1551 129
rect 1500 51 1551 95
rect 1585 161 1639 177
rect 1619 127 1639 161
rect 1585 93 1639 127
rect 1619 59 1639 93
rect 1585 17 1639 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 122 289 156 323
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 494 357 528 391
rect 586 289 620 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 482 391 540 397
rect 482 388 494 391
rect 248 360 494 388
rect 248 357 260 360
rect 202 351 260 357
rect 482 357 494 360
rect 528 357 540 391
rect 482 351 540 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 574 323 632 329
rect 574 320 586 323
rect 156 292 586 320
rect 156 289 168 292
rect 110 283 168 289
rect 574 289 586 292
rect 620 289 632 323
rect 574 283 632 289
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel locali s 310 221 344 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1142 425 1176 459 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1142 85 1176 119 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1230 221 1264 255 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 958 221 992 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1597 221 1631 255 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1505 425 1539 459 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1505 357 1539 391 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1505 85 1539 119 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 dlrbn_2
rlabel metal1 s 0 -48 1656 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1656 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_END 2736830
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2723488
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 41.400 13.600 
<< end >>
