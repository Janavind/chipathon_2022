magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< metal3 >>
rect 10078 1778 14858 2706
<< obsm3 >>
rect 99 1778 4879 2706
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 254 12537
rect 14746 11647 15000 12537
rect 0 11281 15000 11347
rect 0 10625 15000 11221
rect 0 10329 254 10565
rect 14746 10329 15000 10565
rect 0 9673 15000 10269
rect 0 9547 15000 9613
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 7347 254 8037
rect 14746 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 254 6097
rect 14746 5167 15000 6097
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 269 2640 333 2704
rect 351 2640 415 2704
rect 433 2640 497 2704
rect 515 2640 579 2704
rect 597 2640 661 2704
rect 678 2640 742 2704
rect 759 2640 823 2704
rect 840 2640 904 2704
rect 921 2640 985 2704
rect 1002 2640 1066 2704
rect 1083 2640 1147 2704
rect 1164 2640 1228 2704
rect 1245 2640 1309 2704
rect 1326 2640 1390 2704
rect 1407 2640 1471 2704
rect 1488 2640 1552 2704
rect 1569 2640 1633 2704
rect 1650 2640 1714 2704
rect 1731 2640 1795 2704
rect 1812 2640 1876 2704
rect 1893 2640 1957 2704
rect 1974 2640 2038 2704
rect 2055 2640 2119 2704
rect 2136 2640 2200 2704
rect 2217 2640 2281 2704
rect 2298 2640 2362 2704
rect 2379 2640 2443 2704
rect 2460 2640 2524 2704
rect 2541 2640 2605 2704
rect 2622 2640 2686 2704
rect 2703 2640 2767 2704
rect 2784 2640 2848 2704
rect 2865 2640 2929 2704
rect 2946 2640 3010 2704
rect 3027 2640 3091 2704
rect 3108 2640 3172 2704
rect 3189 2640 3253 2704
rect 3270 2640 3334 2704
rect 3351 2640 3415 2704
rect 3432 2640 3496 2704
rect 3513 2640 3577 2704
rect 3594 2640 3658 2704
rect 3675 2640 3739 2704
rect 3756 2640 3820 2704
rect 3837 2640 3901 2704
rect 3918 2640 3982 2704
rect 3999 2640 4063 2704
rect 4080 2640 4144 2704
rect 4161 2640 4225 2704
rect 4242 2640 4306 2704
rect 4323 2640 4387 2704
rect 4404 2640 4468 2704
rect 4485 2640 4549 2704
rect 4566 2640 4630 2704
rect 4647 2640 4711 2704
rect 4728 2640 4792 2704
rect 4809 2640 4873 2704
rect 269 2554 333 2618
rect 351 2554 415 2618
rect 433 2554 497 2618
rect 515 2554 579 2618
rect 597 2554 661 2618
rect 678 2554 742 2618
rect 759 2554 823 2618
rect 840 2554 904 2618
rect 921 2554 985 2618
rect 1002 2554 1066 2618
rect 1083 2554 1147 2618
rect 1164 2554 1228 2618
rect 1245 2554 1309 2618
rect 1326 2554 1390 2618
rect 1407 2554 1471 2618
rect 1488 2554 1552 2618
rect 1569 2554 1633 2618
rect 1650 2554 1714 2618
rect 1731 2554 1795 2618
rect 1812 2554 1876 2618
rect 1893 2554 1957 2618
rect 1974 2554 2038 2618
rect 2055 2554 2119 2618
rect 2136 2554 2200 2618
rect 2217 2554 2281 2618
rect 2298 2554 2362 2618
rect 2379 2554 2443 2618
rect 2460 2554 2524 2618
rect 2541 2554 2605 2618
rect 2622 2554 2686 2618
rect 2703 2554 2767 2618
rect 2784 2554 2848 2618
rect 2865 2554 2929 2618
rect 2946 2554 3010 2618
rect 3027 2554 3091 2618
rect 3108 2554 3172 2618
rect 3189 2554 3253 2618
rect 3270 2554 3334 2618
rect 3351 2554 3415 2618
rect 3432 2554 3496 2618
rect 3513 2554 3577 2618
rect 3594 2554 3658 2618
rect 3675 2554 3739 2618
rect 3756 2554 3820 2618
rect 3837 2554 3901 2618
rect 3918 2554 3982 2618
rect 3999 2554 4063 2618
rect 4080 2554 4144 2618
rect 4161 2554 4225 2618
rect 4242 2554 4306 2618
rect 4323 2554 4387 2618
rect 4404 2554 4468 2618
rect 4485 2554 4549 2618
rect 4566 2554 4630 2618
rect 4647 2554 4711 2618
rect 4728 2554 4792 2618
rect 4809 2554 4873 2618
rect 269 2468 333 2532
rect 351 2468 415 2532
rect 433 2468 497 2532
rect 515 2468 579 2532
rect 597 2468 661 2532
rect 678 2468 742 2532
rect 759 2468 823 2532
rect 840 2468 904 2532
rect 921 2468 985 2532
rect 1002 2468 1066 2532
rect 1083 2468 1147 2532
rect 1164 2468 1228 2532
rect 1245 2468 1309 2532
rect 1326 2468 1390 2532
rect 1407 2468 1471 2532
rect 1488 2468 1552 2532
rect 1569 2468 1633 2532
rect 1650 2468 1714 2532
rect 1731 2468 1795 2532
rect 1812 2468 1876 2532
rect 1893 2468 1957 2532
rect 1974 2468 2038 2532
rect 2055 2468 2119 2532
rect 2136 2468 2200 2532
rect 2217 2468 2281 2532
rect 2298 2468 2362 2532
rect 2379 2468 2443 2532
rect 2460 2468 2524 2532
rect 2541 2468 2605 2532
rect 2622 2468 2686 2532
rect 2703 2468 2767 2532
rect 2784 2468 2848 2532
rect 2865 2468 2929 2532
rect 2946 2468 3010 2532
rect 3027 2468 3091 2532
rect 3108 2468 3172 2532
rect 3189 2468 3253 2532
rect 3270 2468 3334 2532
rect 3351 2468 3415 2532
rect 3432 2468 3496 2532
rect 3513 2468 3577 2532
rect 3594 2468 3658 2532
rect 3675 2468 3739 2532
rect 3756 2468 3820 2532
rect 3837 2468 3901 2532
rect 3918 2468 3982 2532
rect 3999 2468 4063 2532
rect 4080 2468 4144 2532
rect 4161 2468 4225 2532
rect 4242 2468 4306 2532
rect 4323 2468 4387 2532
rect 4404 2468 4468 2532
rect 4485 2468 4549 2532
rect 4566 2468 4630 2532
rect 4647 2468 4711 2532
rect 4728 2468 4792 2532
rect 4809 2468 4873 2532
rect 269 2382 333 2446
rect 351 2382 415 2446
rect 433 2382 497 2446
rect 515 2382 579 2446
rect 597 2382 661 2446
rect 678 2382 742 2446
rect 759 2382 823 2446
rect 840 2382 904 2446
rect 921 2382 985 2446
rect 1002 2382 1066 2446
rect 1083 2382 1147 2446
rect 1164 2382 1228 2446
rect 1245 2382 1309 2446
rect 1326 2382 1390 2446
rect 1407 2382 1471 2446
rect 1488 2382 1552 2446
rect 1569 2382 1633 2446
rect 1650 2382 1714 2446
rect 1731 2382 1795 2446
rect 1812 2382 1876 2446
rect 1893 2382 1957 2446
rect 1974 2382 2038 2446
rect 2055 2382 2119 2446
rect 2136 2382 2200 2446
rect 2217 2382 2281 2446
rect 2298 2382 2362 2446
rect 2379 2382 2443 2446
rect 2460 2382 2524 2446
rect 2541 2382 2605 2446
rect 2622 2382 2686 2446
rect 2703 2382 2767 2446
rect 2784 2382 2848 2446
rect 2865 2382 2929 2446
rect 2946 2382 3010 2446
rect 3027 2382 3091 2446
rect 3108 2382 3172 2446
rect 3189 2382 3253 2446
rect 3270 2382 3334 2446
rect 3351 2382 3415 2446
rect 3432 2382 3496 2446
rect 3513 2382 3577 2446
rect 3594 2382 3658 2446
rect 3675 2382 3739 2446
rect 3756 2382 3820 2446
rect 3837 2382 3901 2446
rect 3918 2382 3982 2446
rect 3999 2382 4063 2446
rect 4080 2382 4144 2446
rect 4161 2382 4225 2446
rect 4242 2382 4306 2446
rect 4323 2382 4387 2446
rect 4404 2382 4468 2446
rect 4485 2382 4549 2446
rect 4566 2382 4630 2446
rect 4647 2382 4711 2446
rect 4728 2382 4792 2446
rect 4809 2382 4873 2446
rect 269 2296 333 2360
rect 351 2296 415 2360
rect 433 2296 497 2360
rect 515 2296 579 2360
rect 597 2296 661 2360
rect 678 2296 742 2360
rect 759 2296 823 2360
rect 840 2296 904 2360
rect 921 2296 985 2360
rect 1002 2296 1066 2360
rect 1083 2296 1147 2360
rect 1164 2296 1228 2360
rect 1245 2296 1309 2360
rect 1326 2296 1390 2360
rect 1407 2296 1471 2360
rect 1488 2296 1552 2360
rect 1569 2296 1633 2360
rect 1650 2296 1714 2360
rect 1731 2296 1795 2360
rect 1812 2296 1876 2360
rect 1893 2296 1957 2360
rect 1974 2296 2038 2360
rect 2055 2296 2119 2360
rect 2136 2296 2200 2360
rect 2217 2296 2281 2360
rect 2298 2296 2362 2360
rect 2379 2296 2443 2360
rect 2460 2296 2524 2360
rect 2541 2296 2605 2360
rect 2622 2296 2686 2360
rect 2703 2296 2767 2360
rect 2784 2296 2848 2360
rect 2865 2296 2929 2360
rect 2946 2296 3010 2360
rect 3027 2296 3091 2360
rect 3108 2296 3172 2360
rect 3189 2296 3253 2360
rect 3270 2296 3334 2360
rect 3351 2296 3415 2360
rect 3432 2296 3496 2360
rect 3513 2296 3577 2360
rect 3594 2296 3658 2360
rect 3675 2296 3739 2360
rect 3756 2296 3820 2360
rect 3837 2296 3901 2360
rect 3918 2296 3982 2360
rect 3999 2296 4063 2360
rect 4080 2296 4144 2360
rect 4161 2296 4225 2360
rect 4242 2296 4306 2360
rect 4323 2296 4387 2360
rect 4404 2296 4468 2360
rect 4485 2296 4549 2360
rect 4566 2296 4630 2360
rect 4647 2296 4711 2360
rect 4728 2296 4792 2360
rect 4809 2296 4873 2360
rect 269 2210 333 2274
rect 351 2210 415 2274
rect 433 2210 497 2274
rect 515 2210 579 2274
rect 597 2210 661 2274
rect 678 2210 742 2274
rect 759 2210 823 2274
rect 840 2210 904 2274
rect 921 2210 985 2274
rect 1002 2210 1066 2274
rect 1083 2210 1147 2274
rect 1164 2210 1228 2274
rect 1245 2210 1309 2274
rect 1326 2210 1390 2274
rect 1407 2210 1471 2274
rect 1488 2210 1552 2274
rect 1569 2210 1633 2274
rect 1650 2210 1714 2274
rect 1731 2210 1795 2274
rect 1812 2210 1876 2274
rect 1893 2210 1957 2274
rect 1974 2210 2038 2274
rect 2055 2210 2119 2274
rect 2136 2210 2200 2274
rect 2217 2210 2281 2274
rect 2298 2210 2362 2274
rect 2379 2210 2443 2274
rect 2460 2210 2524 2274
rect 2541 2210 2605 2274
rect 2622 2210 2686 2274
rect 2703 2210 2767 2274
rect 2784 2210 2848 2274
rect 2865 2210 2929 2274
rect 2946 2210 3010 2274
rect 3027 2210 3091 2274
rect 3108 2210 3172 2274
rect 3189 2210 3253 2274
rect 3270 2210 3334 2274
rect 3351 2210 3415 2274
rect 3432 2210 3496 2274
rect 3513 2210 3577 2274
rect 3594 2210 3658 2274
rect 3675 2210 3739 2274
rect 3756 2210 3820 2274
rect 3837 2210 3901 2274
rect 3918 2210 3982 2274
rect 3999 2210 4063 2274
rect 4080 2210 4144 2274
rect 4161 2210 4225 2274
rect 4242 2210 4306 2274
rect 4323 2210 4387 2274
rect 4404 2210 4468 2274
rect 4485 2210 4549 2274
rect 4566 2210 4630 2274
rect 4647 2210 4711 2274
rect 4728 2210 4792 2274
rect 4809 2210 4873 2274
rect 269 2124 333 2188
rect 351 2124 415 2188
rect 433 2124 497 2188
rect 515 2124 579 2188
rect 597 2124 661 2188
rect 678 2124 742 2188
rect 759 2124 823 2188
rect 840 2124 904 2188
rect 921 2124 985 2188
rect 1002 2124 1066 2188
rect 1083 2124 1147 2188
rect 1164 2124 1228 2188
rect 1245 2124 1309 2188
rect 1326 2124 1390 2188
rect 1407 2124 1471 2188
rect 1488 2124 1552 2188
rect 1569 2124 1633 2188
rect 1650 2124 1714 2188
rect 1731 2124 1795 2188
rect 1812 2124 1876 2188
rect 1893 2124 1957 2188
rect 1974 2124 2038 2188
rect 2055 2124 2119 2188
rect 2136 2124 2200 2188
rect 2217 2124 2281 2188
rect 2298 2124 2362 2188
rect 2379 2124 2443 2188
rect 2460 2124 2524 2188
rect 2541 2124 2605 2188
rect 2622 2124 2686 2188
rect 2703 2124 2767 2188
rect 2784 2124 2848 2188
rect 2865 2124 2929 2188
rect 2946 2124 3010 2188
rect 3027 2124 3091 2188
rect 3108 2124 3172 2188
rect 3189 2124 3253 2188
rect 3270 2124 3334 2188
rect 3351 2124 3415 2188
rect 3432 2124 3496 2188
rect 3513 2124 3577 2188
rect 3594 2124 3658 2188
rect 3675 2124 3739 2188
rect 3756 2124 3820 2188
rect 3837 2124 3901 2188
rect 3918 2124 3982 2188
rect 3999 2124 4063 2188
rect 4080 2124 4144 2188
rect 4161 2124 4225 2188
rect 4242 2124 4306 2188
rect 4323 2124 4387 2188
rect 4404 2124 4468 2188
rect 4485 2124 4549 2188
rect 4566 2124 4630 2188
rect 4647 2124 4711 2188
rect 4728 2124 4792 2188
rect 4809 2124 4873 2188
rect 269 2038 333 2102
rect 351 2038 415 2102
rect 433 2038 497 2102
rect 515 2038 579 2102
rect 597 2038 661 2102
rect 678 2038 742 2102
rect 759 2038 823 2102
rect 840 2038 904 2102
rect 921 2038 985 2102
rect 1002 2038 1066 2102
rect 1083 2038 1147 2102
rect 1164 2038 1228 2102
rect 1245 2038 1309 2102
rect 1326 2038 1390 2102
rect 1407 2038 1471 2102
rect 1488 2038 1552 2102
rect 1569 2038 1633 2102
rect 1650 2038 1714 2102
rect 1731 2038 1795 2102
rect 1812 2038 1876 2102
rect 1893 2038 1957 2102
rect 1974 2038 2038 2102
rect 2055 2038 2119 2102
rect 2136 2038 2200 2102
rect 2217 2038 2281 2102
rect 2298 2038 2362 2102
rect 2379 2038 2443 2102
rect 2460 2038 2524 2102
rect 2541 2038 2605 2102
rect 2622 2038 2686 2102
rect 2703 2038 2767 2102
rect 2784 2038 2848 2102
rect 2865 2038 2929 2102
rect 2946 2038 3010 2102
rect 3027 2038 3091 2102
rect 3108 2038 3172 2102
rect 3189 2038 3253 2102
rect 3270 2038 3334 2102
rect 3351 2038 3415 2102
rect 3432 2038 3496 2102
rect 3513 2038 3577 2102
rect 3594 2038 3658 2102
rect 3675 2038 3739 2102
rect 3756 2038 3820 2102
rect 3837 2038 3901 2102
rect 3918 2038 3982 2102
rect 3999 2038 4063 2102
rect 4080 2038 4144 2102
rect 4161 2038 4225 2102
rect 4242 2038 4306 2102
rect 4323 2038 4387 2102
rect 4404 2038 4468 2102
rect 4485 2038 4549 2102
rect 4566 2038 4630 2102
rect 4647 2038 4711 2102
rect 4728 2038 4792 2102
rect 4809 2038 4873 2102
rect 269 1952 333 2016
rect 351 1952 415 2016
rect 433 1952 497 2016
rect 515 1952 579 2016
rect 597 1952 661 2016
rect 678 1952 742 2016
rect 759 1952 823 2016
rect 840 1952 904 2016
rect 921 1952 985 2016
rect 1002 1952 1066 2016
rect 1083 1952 1147 2016
rect 1164 1952 1228 2016
rect 1245 1952 1309 2016
rect 1326 1952 1390 2016
rect 1407 1952 1471 2016
rect 1488 1952 1552 2016
rect 1569 1952 1633 2016
rect 1650 1952 1714 2016
rect 1731 1952 1795 2016
rect 1812 1952 1876 2016
rect 1893 1952 1957 2016
rect 1974 1952 2038 2016
rect 2055 1952 2119 2016
rect 2136 1952 2200 2016
rect 2217 1952 2281 2016
rect 2298 1952 2362 2016
rect 2379 1952 2443 2016
rect 2460 1952 2524 2016
rect 2541 1952 2605 2016
rect 2622 1952 2686 2016
rect 2703 1952 2767 2016
rect 2784 1952 2848 2016
rect 2865 1952 2929 2016
rect 2946 1952 3010 2016
rect 3027 1952 3091 2016
rect 3108 1952 3172 2016
rect 3189 1952 3253 2016
rect 3270 1952 3334 2016
rect 3351 1952 3415 2016
rect 3432 1952 3496 2016
rect 3513 1952 3577 2016
rect 3594 1952 3658 2016
rect 3675 1952 3739 2016
rect 3756 1952 3820 2016
rect 3837 1952 3901 2016
rect 3918 1952 3982 2016
rect 3999 1952 4063 2016
rect 4080 1952 4144 2016
rect 4161 1952 4225 2016
rect 4242 1952 4306 2016
rect 4323 1952 4387 2016
rect 4404 1952 4468 2016
rect 4485 1952 4549 2016
rect 4566 1952 4630 2016
rect 4647 1952 4711 2016
rect 4728 1952 4792 2016
rect 4809 1952 4873 2016
rect 269 1866 333 1930
rect 351 1866 415 1930
rect 433 1866 497 1930
rect 515 1866 579 1930
rect 597 1866 661 1930
rect 678 1866 742 1930
rect 759 1866 823 1930
rect 840 1866 904 1930
rect 921 1866 985 1930
rect 1002 1866 1066 1930
rect 1083 1866 1147 1930
rect 1164 1866 1228 1930
rect 1245 1866 1309 1930
rect 1326 1866 1390 1930
rect 1407 1866 1471 1930
rect 1488 1866 1552 1930
rect 1569 1866 1633 1930
rect 1650 1866 1714 1930
rect 1731 1866 1795 1930
rect 1812 1866 1876 1930
rect 1893 1866 1957 1930
rect 1974 1866 2038 1930
rect 2055 1866 2119 1930
rect 2136 1866 2200 1930
rect 2217 1866 2281 1930
rect 2298 1866 2362 1930
rect 2379 1866 2443 1930
rect 2460 1866 2524 1930
rect 2541 1866 2605 1930
rect 2622 1866 2686 1930
rect 2703 1866 2767 1930
rect 2784 1866 2848 1930
rect 2865 1866 2929 1930
rect 2946 1866 3010 1930
rect 3027 1866 3091 1930
rect 3108 1866 3172 1930
rect 3189 1866 3253 1930
rect 3270 1866 3334 1930
rect 3351 1866 3415 1930
rect 3432 1866 3496 1930
rect 3513 1866 3577 1930
rect 3594 1866 3658 1930
rect 3675 1866 3739 1930
rect 3756 1866 3820 1930
rect 3837 1866 3901 1930
rect 3918 1866 3982 1930
rect 3999 1866 4063 1930
rect 4080 1866 4144 1930
rect 4161 1866 4225 1930
rect 4242 1866 4306 1930
rect 4323 1866 4387 1930
rect 4404 1866 4468 1930
rect 4485 1866 4549 1930
rect 4566 1866 4630 1930
rect 4647 1866 4711 1930
rect 4728 1866 4792 1930
rect 4809 1866 4873 1930
rect 269 1780 333 1844
rect 351 1780 415 1844
rect 433 1780 497 1844
rect 515 1780 579 1844
rect 597 1780 661 1844
rect 678 1780 742 1844
rect 759 1780 823 1844
rect 840 1780 904 1844
rect 921 1780 985 1844
rect 1002 1780 1066 1844
rect 1083 1780 1147 1844
rect 1164 1780 1228 1844
rect 1245 1780 1309 1844
rect 1326 1780 1390 1844
rect 1407 1780 1471 1844
rect 1488 1780 1552 1844
rect 1569 1780 1633 1844
rect 1650 1780 1714 1844
rect 1731 1780 1795 1844
rect 1812 1780 1876 1844
rect 1893 1780 1957 1844
rect 1974 1780 2038 1844
rect 2055 1780 2119 1844
rect 2136 1780 2200 1844
rect 2217 1780 2281 1844
rect 2298 1780 2362 1844
rect 2379 1780 2443 1844
rect 2460 1780 2524 1844
rect 2541 1780 2605 1844
rect 2622 1780 2686 1844
rect 2703 1780 2767 1844
rect 2784 1780 2848 1844
rect 2865 1780 2929 1844
rect 2946 1780 3010 1844
rect 3027 1780 3091 1844
rect 3108 1780 3172 1844
rect 3189 1780 3253 1844
rect 3270 1780 3334 1844
rect 3351 1780 3415 1844
rect 3432 1780 3496 1844
rect 3513 1780 3577 1844
rect 3594 1780 3658 1844
rect 3675 1780 3739 1844
rect 3756 1780 3820 1844
rect 3837 1780 3901 1844
rect 3918 1780 3982 1844
rect 3999 1780 4063 1844
rect 4080 1780 4144 1844
rect 4161 1780 4225 1844
rect 4242 1780 4306 1844
rect 4323 1780 4387 1844
rect 4404 1780 4468 1844
rect 4485 1780 4549 1844
rect 4566 1780 4630 1844
rect 4647 1780 4711 1844
rect 4728 1780 4792 1844
rect 4809 1780 4873 1844
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< obsm4 >>
rect 334 35077 14666 40000
rect 193 19080 14807 35077
rect 334 13927 14666 19080
rect 193 13787 14807 13927
rect 334 12737 14666 13787
rect 193 12617 14807 12737
rect 334 11567 14666 12617
rect 193 11427 14807 11567
rect 334 10349 14666 10545
rect 193 9327 14807 9467
rect 334 8237 14666 9327
rect 193 8117 14807 8237
rect 334 7267 14666 8117
rect 193 7147 14807 7267
rect 334 6297 14666 7147
rect 193 6177 14807 6297
rect 334 5087 14666 6177
rect 193 4967 14807 5087
rect 334 3877 14666 4967
rect 193 3757 14807 3877
rect 273 2907 14727 3757
rect 193 2787 14807 2907
rect 334 2704 14666 2787
rect 334 2640 351 2704
rect 415 2640 433 2704
rect 497 2640 515 2704
rect 579 2640 597 2704
rect 661 2640 678 2704
rect 742 2640 759 2704
rect 823 2640 840 2704
rect 904 2640 921 2704
rect 985 2640 1002 2704
rect 1066 2640 1083 2704
rect 1147 2640 1164 2704
rect 1228 2640 1245 2704
rect 1309 2640 1326 2704
rect 1390 2640 1407 2704
rect 1471 2640 1488 2704
rect 1552 2640 1569 2704
rect 1633 2640 1650 2704
rect 1714 2640 1731 2704
rect 1795 2640 1812 2704
rect 1876 2640 1893 2704
rect 1957 2640 1974 2704
rect 2038 2640 2055 2704
rect 2119 2640 2136 2704
rect 2200 2640 2217 2704
rect 2281 2640 2298 2704
rect 2362 2640 2379 2704
rect 2443 2640 2460 2704
rect 2524 2640 2541 2704
rect 2605 2640 2622 2704
rect 2686 2640 2703 2704
rect 2767 2640 2784 2704
rect 2848 2640 2865 2704
rect 2929 2640 2946 2704
rect 3010 2640 3027 2704
rect 3091 2640 3108 2704
rect 3172 2640 3189 2704
rect 3253 2640 3270 2704
rect 3334 2640 3351 2704
rect 3415 2640 3432 2704
rect 3496 2640 3513 2704
rect 3577 2640 3594 2704
rect 3658 2640 3675 2704
rect 3739 2640 3756 2704
rect 3820 2640 3837 2704
rect 3901 2640 3918 2704
rect 3982 2640 3999 2704
rect 4063 2640 4080 2704
rect 4144 2640 4161 2704
rect 4225 2640 4242 2704
rect 4306 2640 4323 2704
rect 4387 2640 4404 2704
rect 4468 2640 4485 2704
rect 4549 2640 4566 2704
rect 4630 2640 4647 2704
rect 4711 2640 4728 2704
rect 4792 2640 4809 2704
rect 4873 2640 14666 2704
rect 334 2618 14666 2640
rect 334 2554 351 2618
rect 415 2554 433 2618
rect 497 2554 515 2618
rect 579 2554 597 2618
rect 661 2554 678 2618
rect 742 2554 759 2618
rect 823 2554 840 2618
rect 904 2554 921 2618
rect 985 2554 1002 2618
rect 1066 2554 1083 2618
rect 1147 2554 1164 2618
rect 1228 2554 1245 2618
rect 1309 2554 1326 2618
rect 1390 2554 1407 2618
rect 1471 2554 1488 2618
rect 1552 2554 1569 2618
rect 1633 2554 1650 2618
rect 1714 2554 1731 2618
rect 1795 2554 1812 2618
rect 1876 2554 1893 2618
rect 1957 2554 1974 2618
rect 2038 2554 2055 2618
rect 2119 2554 2136 2618
rect 2200 2554 2217 2618
rect 2281 2554 2298 2618
rect 2362 2554 2379 2618
rect 2443 2554 2460 2618
rect 2524 2554 2541 2618
rect 2605 2554 2622 2618
rect 2686 2554 2703 2618
rect 2767 2554 2784 2618
rect 2848 2554 2865 2618
rect 2929 2554 2946 2618
rect 3010 2554 3027 2618
rect 3091 2554 3108 2618
rect 3172 2554 3189 2618
rect 3253 2554 3270 2618
rect 3334 2554 3351 2618
rect 3415 2554 3432 2618
rect 3496 2554 3513 2618
rect 3577 2554 3594 2618
rect 3658 2554 3675 2618
rect 3739 2554 3756 2618
rect 3820 2554 3837 2618
rect 3901 2554 3918 2618
rect 3982 2554 3999 2618
rect 4063 2554 4080 2618
rect 4144 2554 4161 2618
rect 4225 2554 4242 2618
rect 4306 2554 4323 2618
rect 4387 2554 4404 2618
rect 4468 2554 4485 2618
rect 4549 2554 4566 2618
rect 4630 2554 4647 2618
rect 4711 2554 4728 2618
rect 4792 2554 4809 2618
rect 4873 2554 14666 2618
rect 334 2532 14666 2554
rect 334 2468 351 2532
rect 415 2468 433 2532
rect 497 2468 515 2532
rect 579 2468 597 2532
rect 661 2468 678 2532
rect 742 2468 759 2532
rect 823 2468 840 2532
rect 904 2468 921 2532
rect 985 2468 1002 2532
rect 1066 2468 1083 2532
rect 1147 2468 1164 2532
rect 1228 2468 1245 2532
rect 1309 2468 1326 2532
rect 1390 2468 1407 2532
rect 1471 2468 1488 2532
rect 1552 2468 1569 2532
rect 1633 2468 1650 2532
rect 1714 2468 1731 2532
rect 1795 2468 1812 2532
rect 1876 2468 1893 2532
rect 1957 2468 1974 2532
rect 2038 2468 2055 2532
rect 2119 2468 2136 2532
rect 2200 2468 2217 2532
rect 2281 2468 2298 2532
rect 2362 2468 2379 2532
rect 2443 2468 2460 2532
rect 2524 2468 2541 2532
rect 2605 2468 2622 2532
rect 2686 2468 2703 2532
rect 2767 2468 2784 2532
rect 2848 2468 2865 2532
rect 2929 2468 2946 2532
rect 3010 2468 3027 2532
rect 3091 2468 3108 2532
rect 3172 2468 3189 2532
rect 3253 2468 3270 2532
rect 3334 2468 3351 2532
rect 3415 2468 3432 2532
rect 3496 2468 3513 2532
rect 3577 2468 3594 2532
rect 3658 2468 3675 2532
rect 3739 2468 3756 2532
rect 3820 2468 3837 2532
rect 3901 2468 3918 2532
rect 3982 2468 3999 2532
rect 4063 2468 4080 2532
rect 4144 2468 4161 2532
rect 4225 2468 4242 2532
rect 4306 2468 4323 2532
rect 4387 2468 4404 2532
rect 4468 2468 4485 2532
rect 4549 2468 4566 2532
rect 4630 2468 4647 2532
rect 4711 2468 4728 2532
rect 4792 2468 4809 2532
rect 4873 2468 14666 2532
rect 334 2446 14666 2468
rect 334 2382 351 2446
rect 415 2382 433 2446
rect 497 2382 515 2446
rect 579 2382 597 2446
rect 661 2382 678 2446
rect 742 2382 759 2446
rect 823 2382 840 2446
rect 904 2382 921 2446
rect 985 2382 1002 2446
rect 1066 2382 1083 2446
rect 1147 2382 1164 2446
rect 1228 2382 1245 2446
rect 1309 2382 1326 2446
rect 1390 2382 1407 2446
rect 1471 2382 1488 2446
rect 1552 2382 1569 2446
rect 1633 2382 1650 2446
rect 1714 2382 1731 2446
rect 1795 2382 1812 2446
rect 1876 2382 1893 2446
rect 1957 2382 1974 2446
rect 2038 2382 2055 2446
rect 2119 2382 2136 2446
rect 2200 2382 2217 2446
rect 2281 2382 2298 2446
rect 2362 2382 2379 2446
rect 2443 2382 2460 2446
rect 2524 2382 2541 2446
rect 2605 2382 2622 2446
rect 2686 2382 2703 2446
rect 2767 2382 2784 2446
rect 2848 2382 2865 2446
rect 2929 2382 2946 2446
rect 3010 2382 3027 2446
rect 3091 2382 3108 2446
rect 3172 2382 3189 2446
rect 3253 2382 3270 2446
rect 3334 2382 3351 2446
rect 3415 2382 3432 2446
rect 3496 2382 3513 2446
rect 3577 2382 3594 2446
rect 3658 2382 3675 2446
rect 3739 2382 3756 2446
rect 3820 2382 3837 2446
rect 3901 2382 3918 2446
rect 3982 2382 3999 2446
rect 4063 2382 4080 2446
rect 4144 2382 4161 2446
rect 4225 2382 4242 2446
rect 4306 2382 4323 2446
rect 4387 2382 4404 2446
rect 4468 2382 4485 2446
rect 4549 2382 4566 2446
rect 4630 2382 4647 2446
rect 4711 2382 4728 2446
rect 4792 2382 4809 2446
rect 4873 2382 14666 2446
rect 334 2360 14666 2382
rect 334 2296 351 2360
rect 415 2296 433 2360
rect 497 2296 515 2360
rect 579 2296 597 2360
rect 661 2296 678 2360
rect 742 2296 759 2360
rect 823 2296 840 2360
rect 904 2296 921 2360
rect 985 2296 1002 2360
rect 1066 2296 1083 2360
rect 1147 2296 1164 2360
rect 1228 2296 1245 2360
rect 1309 2296 1326 2360
rect 1390 2296 1407 2360
rect 1471 2296 1488 2360
rect 1552 2296 1569 2360
rect 1633 2296 1650 2360
rect 1714 2296 1731 2360
rect 1795 2296 1812 2360
rect 1876 2296 1893 2360
rect 1957 2296 1974 2360
rect 2038 2296 2055 2360
rect 2119 2296 2136 2360
rect 2200 2296 2217 2360
rect 2281 2296 2298 2360
rect 2362 2296 2379 2360
rect 2443 2296 2460 2360
rect 2524 2296 2541 2360
rect 2605 2296 2622 2360
rect 2686 2296 2703 2360
rect 2767 2296 2784 2360
rect 2848 2296 2865 2360
rect 2929 2296 2946 2360
rect 3010 2296 3027 2360
rect 3091 2296 3108 2360
rect 3172 2296 3189 2360
rect 3253 2296 3270 2360
rect 3334 2296 3351 2360
rect 3415 2296 3432 2360
rect 3496 2296 3513 2360
rect 3577 2296 3594 2360
rect 3658 2296 3675 2360
rect 3739 2296 3756 2360
rect 3820 2296 3837 2360
rect 3901 2296 3918 2360
rect 3982 2296 3999 2360
rect 4063 2296 4080 2360
rect 4144 2296 4161 2360
rect 4225 2296 4242 2360
rect 4306 2296 4323 2360
rect 4387 2296 4404 2360
rect 4468 2296 4485 2360
rect 4549 2296 4566 2360
rect 4630 2296 4647 2360
rect 4711 2296 4728 2360
rect 4792 2296 4809 2360
rect 4873 2296 14666 2360
rect 334 2274 14666 2296
rect 334 2210 351 2274
rect 415 2210 433 2274
rect 497 2210 515 2274
rect 579 2210 597 2274
rect 661 2210 678 2274
rect 742 2210 759 2274
rect 823 2210 840 2274
rect 904 2210 921 2274
rect 985 2210 1002 2274
rect 1066 2210 1083 2274
rect 1147 2210 1164 2274
rect 1228 2210 1245 2274
rect 1309 2210 1326 2274
rect 1390 2210 1407 2274
rect 1471 2210 1488 2274
rect 1552 2210 1569 2274
rect 1633 2210 1650 2274
rect 1714 2210 1731 2274
rect 1795 2210 1812 2274
rect 1876 2210 1893 2274
rect 1957 2210 1974 2274
rect 2038 2210 2055 2274
rect 2119 2210 2136 2274
rect 2200 2210 2217 2274
rect 2281 2210 2298 2274
rect 2362 2210 2379 2274
rect 2443 2210 2460 2274
rect 2524 2210 2541 2274
rect 2605 2210 2622 2274
rect 2686 2210 2703 2274
rect 2767 2210 2784 2274
rect 2848 2210 2865 2274
rect 2929 2210 2946 2274
rect 3010 2210 3027 2274
rect 3091 2210 3108 2274
rect 3172 2210 3189 2274
rect 3253 2210 3270 2274
rect 3334 2210 3351 2274
rect 3415 2210 3432 2274
rect 3496 2210 3513 2274
rect 3577 2210 3594 2274
rect 3658 2210 3675 2274
rect 3739 2210 3756 2274
rect 3820 2210 3837 2274
rect 3901 2210 3918 2274
rect 3982 2210 3999 2274
rect 4063 2210 4080 2274
rect 4144 2210 4161 2274
rect 4225 2210 4242 2274
rect 4306 2210 4323 2274
rect 4387 2210 4404 2274
rect 4468 2210 4485 2274
rect 4549 2210 4566 2274
rect 4630 2210 4647 2274
rect 4711 2210 4728 2274
rect 4792 2210 4809 2274
rect 4873 2210 14666 2274
rect 334 2188 14666 2210
rect 334 2124 351 2188
rect 415 2124 433 2188
rect 497 2124 515 2188
rect 579 2124 597 2188
rect 661 2124 678 2188
rect 742 2124 759 2188
rect 823 2124 840 2188
rect 904 2124 921 2188
rect 985 2124 1002 2188
rect 1066 2124 1083 2188
rect 1147 2124 1164 2188
rect 1228 2124 1245 2188
rect 1309 2124 1326 2188
rect 1390 2124 1407 2188
rect 1471 2124 1488 2188
rect 1552 2124 1569 2188
rect 1633 2124 1650 2188
rect 1714 2124 1731 2188
rect 1795 2124 1812 2188
rect 1876 2124 1893 2188
rect 1957 2124 1974 2188
rect 2038 2124 2055 2188
rect 2119 2124 2136 2188
rect 2200 2124 2217 2188
rect 2281 2124 2298 2188
rect 2362 2124 2379 2188
rect 2443 2124 2460 2188
rect 2524 2124 2541 2188
rect 2605 2124 2622 2188
rect 2686 2124 2703 2188
rect 2767 2124 2784 2188
rect 2848 2124 2865 2188
rect 2929 2124 2946 2188
rect 3010 2124 3027 2188
rect 3091 2124 3108 2188
rect 3172 2124 3189 2188
rect 3253 2124 3270 2188
rect 3334 2124 3351 2188
rect 3415 2124 3432 2188
rect 3496 2124 3513 2188
rect 3577 2124 3594 2188
rect 3658 2124 3675 2188
rect 3739 2124 3756 2188
rect 3820 2124 3837 2188
rect 3901 2124 3918 2188
rect 3982 2124 3999 2188
rect 4063 2124 4080 2188
rect 4144 2124 4161 2188
rect 4225 2124 4242 2188
rect 4306 2124 4323 2188
rect 4387 2124 4404 2188
rect 4468 2124 4485 2188
rect 4549 2124 4566 2188
rect 4630 2124 4647 2188
rect 4711 2124 4728 2188
rect 4792 2124 4809 2188
rect 4873 2124 14666 2188
rect 334 2102 14666 2124
rect 334 2038 351 2102
rect 415 2038 433 2102
rect 497 2038 515 2102
rect 579 2038 597 2102
rect 661 2038 678 2102
rect 742 2038 759 2102
rect 823 2038 840 2102
rect 904 2038 921 2102
rect 985 2038 1002 2102
rect 1066 2038 1083 2102
rect 1147 2038 1164 2102
rect 1228 2038 1245 2102
rect 1309 2038 1326 2102
rect 1390 2038 1407 2102
rect 1471 2038 1488 2102
rect 1552 2038 1569 2102
rect 1633 2038 1650 2102
rect 1714 2038 1731 2102
rect 1795 2038 1812 2102
rect 1876 2038 1893 2102
rect 1957 2038 1974 2102
rect 2038 2038 2055 2102
rect 2119 2038 2136 2102
rect 2200 2038 2217 2102
rect 2281 2038 2298 2102
rect 2362 2038 2379 2102
rect 2443 2038 2460 2102
rect 2524 2038 2541 2102
rect 2605 2038 2622 2102
rect 2686 2038 2703 2102
rect 2767 2038 2784 2102
rect 2848 2038 2865 2102
rect 2929 2038 2946 2102
rect 3010 2038 3027 2102
rect 3091 2038 3108 2102
rect 3172 2038 3189 2102
rect 3253 2038 3270 2102
rect 3334 2038 3351 2102
rect 3415 2038 3432 2102
rect 3496 2038 3513 2102
rect 3577 2038 3594 2102
rect 3658 2038 3675 2102
rect 3739 2038 3756 2102
rect 3820 2038 3837 2102
rect 3901 2038 3918 2102
rect 3982 2038 3999 2102
rect 4063 2038 4080 2102
rect 4144 2038 4161 2102
rect 4225 2038 4242 2102
rect 4306 2038 4323 2102
rect 4387 2038 4404 2102
rect 4468 2038 4485 2102
rect 4549 2038 4566 2102
rect 4630 2038 4647 2102
rect 4711 2038 4728 2102
rect 4792 2038 4809 2102
rect 4873 2038 14666 2102
rect 334 2016 14666 2038
rect 334 1952 351 2016
rect 415 1952 433 2016
rect 497 1952 515 2016
rect 579 1952 597 2016
rect 661 1952 678 2016
rect 742 1952 759 2016
rect 823 1952 840 2016
rect 904 1952 921 2016
rect 985 1952 1002 2016
rect 1066 1952 1083 2016
rect 1147 1952 1164 2016
rect 1228 1952 1245 2016
rect 1309 1952 1326 2016
rect 1390 1952 1407 2016
rect 1471 1952 1488 2016
rect 1552 1952 1569 2016
rect 1633 1952 1650 2016
rect 1714 1952 1731 2016
rect 1795 1952 1812 2016
rect 1876 1952 1893 2016
rect 1957 1952 1974 2016
rect 2038 1952 2055 2016
rect 2119 1952 2136 2016
rect 2200 1952 2217 2016
rect 2281 1952 2298 2016
rect 2362 1952 2379 2016
rect 2443 1952 2460 2016
rect 2524 1952 2541 2016
rect 2605 1952 2622 2016
rect 2686 1952 2703 2016
rect 2767 1952 2784 2016
rect 2848 1952 2865 2016
rect 2929 1952 2946 2016
rect 3010 1952 3027 2016
rect 3091 1952 3108 2016
rect 3172 1952 3189 2016
rect 3253 1952 3270 2016
rect 3334 1952 3351 2016
rect 3415 1952 3432 2016
rect 3496 1952 3513 2016
rect 3577 1952 3594 2016
rect 3658 1952 3675 2016
rect 3739 1952 3756 2016
rect 3820 1952 3837 2016
rect 3901 1952 3918 2016
rect 3982 1952 3999 2016
rect 4063 1952 4080 2016
rect 4144 1952 4161 2016
rect 4225 1952 4242 2016
rect 4306 1952 4323 2016
rect 4387 1952 4404 2016
rect 4468 1952 4485 2016
rect 4549 1952 4566 2016
rect 4630 1952 4647 2016
rect 4711 1952 4728 2016
rect 4792 1952 4809 2016
rect 4873 1952 14666 2016
rect 334 1930 14666 1952
rect 334 1866 351 1930
rect 415 1866 433 1930
rect 497 1866 515 1930
rect 579 1866 597 1930
rect 661 1866 678 1930
rect 742 1866 759 1930
rect 823 1866 840 1930
rect 904 1866 921 1930
rect 985 1866 1002 1930
rect 1066 1866 1083 1930
rect 1147 1866 1164 1930
rect 1228 1866 1245 1930
rect 1309 1866 1326 1930
rect 1390 1866 1407 1930
rect 1471 1866 1488 1930
rect 1552 1866 1569 1930
rect 1633 1866 1650 1930
rect 1714 1866 1731 1930
rect 1795 1866 1812 1930
rect 1876 1866 1893 1930
rect 1957 1866 1974 1930
rect 2038 1866 2055 1930
rect 2119 1866 2136 1930
rect 2200 1866 2217 1930
rect 2281 1866 2298 1930
rect 2362 1866 2379 1930
rect 2443 1866 2460 1930
rect 2524 1866 2541 1930
rect 2605 1866 2622 1930
rect 2686 1866 2703 1930
rect 2767 1866 2784 1930
rect 2848 1866 2865 1930
rect 2929 1866 2946 1930
rect 3010 1866 3027 1930
rect 3091 1866 3108 1930
rect 3172 1866 3189 1930
rect 3253 1866 3270 1930
rect 3334 1866 3351 1930
rect 3415 1866 3432 1930
rect 3496 1866 3513 1930
rect 3577 1866 3594 1930
rect 3658 1866 3675 1930
rect 3739 1866 3756 1930
rect 3820 1866 3837 1930
rect 3901 1866 3918 1930
rect 3982 1866 3999 1930
rect 4063 1866 4080 1930
rect 4144 1866 4161 1930
rect 4225 1866 4242 1930
rect 4306 1866 4323 1930
rect 4387 1866 4404 1930
rect 4468 1866 4485 1930
rect 4549 1866 4566 1930
rect 4630 1866 4647 1930
rect 4711 1866 4728 1930
rect 4792 1866 4809 1930
rect 4873 1866 14666 1930
rect 334 1844 14666 1866
rect 334 1780 351 1844
rect 415 1780 433 1844
rect 497 1780 515 1844
rect 579 1780 597 1844
rect 661 1780 678 1844
rect 742 1780 759 1844
rect 823 1780 840 1844
rect 904 1780 921 1844
rect 985 1780 1002 1844
rect 1066 1780 1083 1844
rect 1147 1780 1164 1844
rect 1228 1780 1245 1844
rect 1309 1780 1326 1844
rect 1390 1780 1407 1844
rect 1471 1780 1488 1844
rect 1552 1780 1569 1844
rect 1633 1780 1650 1844
rect 1714 1780 1731 1844
rect 1795 1780 1812 1844
rect 1876 1780 1893 1844
rect 1957 1780 1974 1844
rect 2038 1780 2055 1844
rect 2119 1780 2136 1844
rect 2200 1780 2217 1844
rect 2281 1780 2298 1844
rect 2362 1780 2379 1844
rect 2443 1780 2460 1844
rect 2524 1780 2541 1844
rect 2605 1780 2622 1844
rect 2686 1780 2703 1844
rect 2767 1780 2784 1844
rect 2848 1780 2865 1844
rect 2929 1780 2946 1844
rect 3010 1780 3027 1844
rect 3091 1780 3108 1844
rect 3172 1780 3189 1844
rect 3253 1780 3270 1844
rect 3334 1780 3351 1844
rect 3415 1780 3432 1844
rect 3496 1780 3513 1844
rect 3577 1780 3594 1844
rect 3658 1780 3675 1844
rect 3739 1780 3756 1844
rect 3820 1780 3837 1844
rect 3901 1780 3918 1844
rect 3982 1780 3999 1844
rect 4063 1780 4080 1844
rect 4144 1780 4161 1844
rect 4225 1780 4242 1844
rect 4306 1780 4323 1844
rect 4387 1780 4404 1844
rect 4468 1780 4485 1844
rect 4549 1780 4566 1844
rect 4630 1780 4647 1844
rect 4711 1780 4728 1844
rect 4792 1780 4809 1844
rect 4873 1780 14666 1844
rect 334 1697 14666 1780
rect 193 1577 14807 1697
rect 334 407 14666 1577
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 18997
rect 0 12837 254 13687
rect 0 11667 254 12517
rect 0 9547 254 11347
rect 0 8337 254 9227
rect 0 7368 254 8017
rect 14746 14007 15000 18997
rect 14746 12837 15000 13687
rect 14746 11667 15000 12517
rect 14746 9547 15000 11347
rect 14746 8337 15000 9227
rect 14746 7368 15000 8017
rect 0 6397 254 7047
rect 0 5187 254 6077
rect 0 3977 254 4867
rect 14746 6397 15000 7047
rect 14746 5187 15000 6077
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 0 427 254 1477
rect 14746 1797 15000 2687
rect 14746 427 15000 1477
<< obsm5 >>
rect 574 34837 14426 40000
rect 0 19317 15000 34837
rect 574 7368 14426 19317
rect 0 7367 15000 7368
rect 574 3657 14426 7367
rect 513 3007 14487 3657
rect 574 427 14426 3007
<< labels >>
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 1 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 1 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 1 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 1 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 1 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 1 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 1 nsew power bidirectional
rlabel metal4 s 0 3957 254 4887 6 VDDIO
port 1 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 2 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 2 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 2 nsew power bidirectional
rlabel metal4 s 0 407 254 1497 6 VCCHIB
port 2 nsew power bidirectional
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9547 15000 9613 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 7347 254 8037 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 11281 15000 11347 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 4 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 4 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 4 nsew power bidirectional
rlabel metal4 s 0 12817 254 13707 6 VDDIO_Q
port 4 nsew power bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 5 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 5 nsew ground bidirectional
rlabel metal4 s 0 11647 254 12537 6 VSSIO_Q
port 5 nsew ground bidirectional
rlabel metal4 s 14746 11647 15000 12537 6 VSSIO_Q
port 5 nsew ground bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal4 s 0 6377 254 7067 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal4 s 0 35157 254 40000 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 8 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 0 1777 254 2707 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10078 1778 14858 2706 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14800 2652 14840 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14800 2566 14840 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14800 2480 14840 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14800 2394 14840 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14800 2308 14840 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14800 2222 14840 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14800 2136 14840 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14800 2050 14840 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14800 1964 14840 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14800 1878 14840 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14800 1792 14840 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14719 2652 14759 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14719 2566 14759 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14719 2480 14759 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14719 2394 14759 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14719 2308 14759 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14719 2222 14759 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14719 2136 14759 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14719 2050 14759 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14719 1964 14759 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14719 1878 14759 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14719 1792 14759 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14638 2652 14678 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14638 2566 14678 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14638 2480 14678 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14638 2394 14678 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14638 2308 14678 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14638 2222 14678 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14638 2136 14678 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14638 2050 14678 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14638 1964 14678 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14638 1878 14678 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14638 1792 14678 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14557 2652 14597 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14557 2566 14597 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14557 2480 14597 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14557 2394 14597 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14557 2308 14597 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14557 2222 14597 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14557 2136 14597 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14557 2050 14597 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14557 1964 14597 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14557 1878 14597 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14557 1792 14597 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14476 2652 14516 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14476 2566 14516 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14476 2480 14516 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14476 2394 14516 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14476 2308 14516 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14476 2222 14516 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14476 2136 14516 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14476 2050 14516 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14476 1964 14516 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14476 1878 14516 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14476 1792 14516 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14395 2652 14435 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14395 2566 14435 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14395 2480 14435 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14395 2394 14435 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14395 2308 14435 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14395 2222 14435 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14395 2136 14435 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14395 2050 14435 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14395 1964 14435 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14395 1878 14435 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14395 1792 14435 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14314 2652 14354 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14314 2566 14354 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14314 2480 14354 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14314 2394 14354 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14314 2308 14354 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14314 2222 14354 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14314 2136 14354 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14314 2050 14354 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14314 1964 14354 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14314 1878 14354 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14314 1792 14354 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14233 2652 14273 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14233 2566 14273 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14233 2480 14273 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14233 2394 14273 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14233 2308 14273 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14233 2222 14273 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14233 2136 14273 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14233 2050 14273 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14233 1964 14273 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14233 1878 14273 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14233 1792 14273 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14152 2652 14192 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14152 2566 14192 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14152 2480 14192 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14152 2394 14192 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14152 2308 14192 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14152 2222 14192 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14152 2136 14192 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14152 2050 14192 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14152 1964 14192 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14152 1878 14192 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14152 1792 14192 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14071 2652 14111 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14071 2566 14111 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14071 2480 14111 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14071 2394 14111 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14071 2308 14111 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14071 2222 14111 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14071 2136 14111 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14071 2050 14111 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14071 1964 14111 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14071 1878 14111 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 14071 1792 14111 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13990 2652 14030 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13990 2566 14030 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13990 2480 14030 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13990 2394 14030 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13990 2308 14030 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13990 2222 14030 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13990 2136 14030 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13990 2050 14030 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13990 1964 14030 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13990 1878 14030 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13990 1792 14030 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13909 2652 13949 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13909 2566 13949 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13909 2480 13949 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13909 2394 13949 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13909 2308 13949 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13909 2222 13949 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13909 2136 13949 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13909 2050 13949 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13909 1964 13949 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13909 1878 13949 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13909 1792 13949 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13828 2652 13868 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13828 2566 13868 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13828 2480 13868 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13828 2394 13868 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13828 2308 13868 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13828 2222 13868 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13828 2136 13868 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13828 2050 13868 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13828 1964 13868 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13828 1878 13868 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13828 1792 13868 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13747 2652 13787 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13747 2566 13787 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13747 2480 13787 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13747 2394 13787 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13747 2308 13787 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13747 2222 13787 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13747 2136 13787 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13747 2050 13787 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13747 1964 13787 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13747 1878 13787 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13747 1792 13787 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13666 2652 13706 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13666 2566 13706 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13666 2480 13706 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13666 2394 13706 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13666 2308 13706 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13666 2222 13706 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13666 2136 13706 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13666 2050 13706 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13666 1964 13706 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13666 1878 13706 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13666 1792 13706 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13585 2652 13625 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13585 2566 13625 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13585 2480 13625 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13585 2394 13625 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13585 2308 13625 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13585 2222 13625 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13585 2136 13625 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13585 2050 13625 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13585 1964 13625 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13585 1878 13625 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13585 1792 13625 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13504 2652 13544 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13504 2566 13544 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13504 2480 13544 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13504 2394 13544 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13504 2308 13544 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13504 2222 13544 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13504 2136 13544 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13504 2050 13544 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13504 1964 13544 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13504 1878 13544 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13504 1792 13544 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13423 2652 13463 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13423 2566 13463 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13423 2480 13463 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13423 2394 13463 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13423 2308 13463 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13423 2222 13463 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13423 2136 13463 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13423 2050 13463 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13423 1964 13463 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13423 1878 13463 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13423 1792 13463 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13342 2652 13382 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13342 2566 13382 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13342 2480 13382 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13342 2394 13382 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13342 2308 13382 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13342 2222 13382 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13342 2136 13382 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13342 2050 13382 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13342 1964 13382 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13342 1878 13382 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13342 1792 13382 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13261 2652 13301 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13261 2566 13301 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13261 2480 13301 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13261 2394 13301 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13261 2308 13301 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13261 2222 13301 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13261 2136 13301 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13261 2050 13301 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13261 1964 13301 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13261 1878 13301 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13261 1792 13301 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13180 2652 13220 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13180 2566 13220 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13180 2480 13220 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13180 2394 13220 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13180 2308 13220 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13180 2222 13220 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13180 2136 13220 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13180 2050 13220 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13180 1964 13220 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13180 1878 13220 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13180 1792 13220 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13099 2652 13139 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13099 2566 13139 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13099 2480 13139 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13099 2394 13139 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13099 2308 13139 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13099 2222 13139 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13099 2136 13139 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13099 2050 13139 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13099 1964 13139 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13099 1878 13139 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13099 1792 13139 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13018 2652 13058 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13018 2566 13058 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13018 2480 13058 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13018 2394 13058 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13018 2308 13058 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13018 2222 13058 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13018 2136 13058 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13018 2050 13058 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13018 1964 13058 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13018 1878 13058 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 13018 1792 13058 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12937 2652 12977 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12937 2566 12977 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12937 2480 12977 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12937 2394 12977 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12937 2308 12977 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12937 2222 12977 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12937 2136 12977 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12937 2050 12977 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12937 1964 12977 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12937 1878 12977 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12937 1792 12977 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12856 2652 12896 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12856 2566 12896 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12856 2480 12896 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12856 2394 12896 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12856 2308 12896 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12856 2222 12896 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12856 2136 12896 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12856 2050 12896 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12856 1964 12896 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12856 1878 12896 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12856 1792 12896 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12775 2652 12815 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12775 2566 12815 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12775 2480 12815 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12775 2394 12815 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12775 2308 12815 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12775 2222 12815 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12775 2136 12815 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12775 2050 12815 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12775 1964 12815 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12775 1878 12815 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12775 1792 12815 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12694 2652 12734 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12694 2566 12734 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12694 2480 12734 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12694 2394 12734 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12694 2308 12734 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12694 2222 12734 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12694 2136 12734 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12694 2050 12734 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12694 1964 12734 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12694 1878 12734 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12694 1792 12734 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12613 2652 12653 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12613 2566 12653 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12613 2480 12653 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12613 2394 12653 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12613 2308 12653 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12613 2222 12653 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12613 2136 12653 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12613 2050 12653 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12613 1964 12653 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12613 1878 12653 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12613 1792 12653 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12532 2652 12572 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12532 2566 12572 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12532 2480 12572 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12532 2394 12572 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12532 2308 12572 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12532 2222 12572 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12532 2136 12572 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12532 2050 12572 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12532 1964 12572 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12532 1878 12572 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12532 1792 12572 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12451 2652 12491 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12451 2566 12491 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12451 2480 12491 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12451 2394 12491 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12451 2308 12491 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12451 2222 12491 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12451 2136 12491 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12451 2050 12491 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12451 1964 12491 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12451 1878 12491 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12451 1792 12491 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12370 2652 12410 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12370 2566 12410 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12370 2480 12410 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12370 2394 12410 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12370 2308 12410 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12370 2222 12410 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12370 2136 12410 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12370 2050 12410 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12370 1964 12410 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12370 1878 12410 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12370 1792 12410 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12289 2652 12329 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12289 2566 12329 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12289 2480 12329 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12289 2394 12329 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12289 2308 12329 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12289 2222 12329 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12289 2136 12329 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12289 2050 12329 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12289 1964 12329 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12289 1878 12329 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12289 1792 12329 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12208 2652 12248 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12208 2566 12248 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12208 2480 12248 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12208 2394 12248 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12208 2308 12248 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12208 2222 12248 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12208 2136 12248 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12208 2050 12248 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12208 1964 12248 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12208 1878 12248 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12208 1792 12248 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12127 2652 12167 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12127 2566 12167 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12127 2480 12167 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12127 2394 12167 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12127 2308 12167 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12127 2222 12167 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12127 2136 12167 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12127 2050 12167 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12127 1964 12167 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12127 1878 12167 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12127 1792 12167 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12046 2652 12086 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12046 2566 12086 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12046 2480 12086 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12046 2394 12086 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12046 2308 12086 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12046 2222 12086 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12046 2136 12086 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12046 2050 12086 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12046 1964 12086 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12046 1878 12086 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 12046 1792 12086 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11965 2652 12005 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11965 2566 12005 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11965 2480 12005 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11965 2394 12005 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11965 2308 12005 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11965 2222 12005 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11965 2136 12005 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11965 2050 12005 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11965 1964 12005 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11965 1878 12005 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11965 1792 12005 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11884 2652 11924 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11884 2566 11924 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11884 2480 11924 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11884 2394 11924 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11884 2308 11924 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11884 2222 11924 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11884 2136 11924 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11884 2050 11924 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11884 1964 11924 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11884 1878 11924 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11884 1792 11924 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11803 2652 11843 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11803 2566 11843 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11803 2480 11843 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11803 2394 11843 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11803 2308 11843 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11803 2222 11843 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11803 2136 11843 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11803 2050 11843 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11803 1964 11843 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11803 1878 11843 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11803 1792 11843 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11722 2652 11762 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11722 2566 11762 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11722 2480 11762 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11722 2394 11762 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11722 2308 11762 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11722 2222 11762 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11722 2136 11762 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11722 2050 11762 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11722 1964 11762 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11722 1878 11762 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11722 1792 11762 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11641 2652 11681 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11641 2566 11681 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11641 2480 11681 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11641 2394 11681 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11641 2308 11681 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11641 2222 11681 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11641 2136 11681 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11641 2050 11681 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11641 1964 11681 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11641 1878 11681 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11641 1792 11681 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11560 2652 11600 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11560 2566 11600 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11560 2480 11600 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11560 2394 11600 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11560 2308 11600 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11560 2222 11600 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11560 2136 11600 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11560 2050 11600 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11560 1964 11600 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11560 1878 11600 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11560 1792 11600 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11479 2652 11519 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11479 2566 11519 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11479 2480 11519 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11479 2394 11519 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11479 2308 11519 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11479 2222 11519 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11479 2136 11519 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11479 2050 11519 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11479 1964 11519 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11479 1878 11519 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11479 1792 11519 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11398 2652 11438 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11398 2566 11438 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11398 2480 11438 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11398 2394 11438 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11398 2308 11438 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11398 2222 11438 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11398 2136 11438 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11398 2050 11438 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11398 1964 11438 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11398 1878 11438 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11398 1792 11438 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11317 2652 11357 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11317 2566 11357 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11317 2480 11357 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11317 2394 11357 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11317 2308 11357 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11317 2222 11357 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11317 2136 11357 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11317 2050 11357 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11317 1964 11357 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11317 1878 11357 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11317 1792 11357 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11236 2652 11276 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11236 2566 11276 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11236 2480 11276 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11236 2394 11276 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11236 2308 11276 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11236 2222 11276 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11236 2136 11276 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11236 2050 11276 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11236 1964 11276 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11236 1878 11276 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11236 1792 11276 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11155 2652 11195 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11155 2566 11195 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11155 2480 11195 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11155 2394 11195 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11155 2308 11195 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11155 2222 11195 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11155 2136 11195 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11155 2050 11195 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11155 1964 11195 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11155 1878 11195 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11155 1792 11195 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11074 2652 11114 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11074 2566 11114 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11074 2480 11114 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11074 2394 11114 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11074 2308 11114 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11074 2222 11114 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11074 2136 11114 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11074 2050 11114 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11074 1964 11114 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11074 1878 11114 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 11074 1792 11114 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10993 2652 11033 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10993 2566 11033 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10993 2480 11033 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10993 2394 11033 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10993 2308 11033 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10993 2222 11033 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10993 2136 11033 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10993 2050 11033 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10993 1964 11033 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10993 1878 11033 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10993 1792 11033 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10912 2652 10952 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10912 2566 10952 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10912 2480 10952 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10912 2394 10952 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10912 2308 10952 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10912 2222 10952 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10912 2136 10952 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10912 2050 10952 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10912 1964 10952 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10912 1878 10952 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10912 1792 10952 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10831 2652 10871 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10831 2566 10871 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10831 2480 10871 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10831 2394 10871 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10831 2308 10871 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10831 2222 10871 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10831 2136 10871 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10831 2050 10871 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10831 1964 10871 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10831 1878 10871 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10831 1792 10871 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10750 2652 10790 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10750 2566 10790 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10750 2480 10790 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10750 2394 10790 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10750 2308 10790 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10750 2222 10790 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10750 2136 10790 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10750 2050 10790 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10750 1964 10790 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10750 1878 10790 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10750 1792 10790 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10669 2652 10709 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10669 2566 10709 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10669 2480 10709 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10669 2394 10709 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10669 2308 10709 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10669 2222 10709 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10669 2136 10709 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10669 2050 10709 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10669 1964 10709 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10669 1878 10709 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10669 1792 10709 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10588 2652 10628 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10588 2566 10628 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10588 2480 10628 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10588 2394 10628 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10588 2308 10628 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10588 2222 10628 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10588 2136 10628 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10588 2050 10628 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10588 1964 10628 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10588 1878 10628 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10588 1792 10628 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10506 2652 10546 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10506 2566 10546 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10506 2480 10546 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10506 2394 10546 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10506 2308 10546 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10506 2222 10546 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10506 2136 10546 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10506 2050 10546 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10506 1964 10546 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10506 1878 10546 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10506 1792 10546 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10424 2652 10464 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10424 2566 10464 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10424 2480 10464 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10424 2394 10464 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10424 2308 10464 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10424 2222 10464 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10424 2136 10464 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10424 2050 10464 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10424 1964 10464 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10424 1878 10464 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10424 1792 10464 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10342 2652 10382 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10342 2566 10382 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10342 2480 10382 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10342 2394 10382 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10342 2308 10382 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10342 2222 10382 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10342 2136 10382 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10342 2050 10382 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10342 1964 10382 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10342 1878 10382 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10342 1792 10382 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10260 2652 10300 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10260 2566 10300 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10260 2480 10300 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10260 2394 10300 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10260 2308 10300 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10260 2222 10300 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10260 2136 10300 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10260 2050 10300 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10260 1964 10300 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10260 1878 10300 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10260 1792 10300 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10178 2652 10218 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10178 2566 10218 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10178 2480 10218 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10178 2394 10218 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10178 2308 10218 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10178 2222 10218 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10178 2136 10218 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10178 2050 10218 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10178 1964 10218 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10178 1878 10218 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10178 1792 10218 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10096 2652 10136 2692 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10096 2566 10136 2606 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10096 2480 10136 2520 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10096 2394 10136 2434 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10096 2308 10136 2348 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10096 2222 10136 2262 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10096 2136 10136 2176 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10096 2050 10136 2090 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10096 1964 10136 2004 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10096 1878 10136 1918 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 10096 1792 10136 1832 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4809 2640 4873 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4809 2640 4873 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4809 2554 4873 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4809 2554 4873 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4809 2468 4873 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4809 2468 4873 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4809 2382 4873 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4809 2382 4873 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4809 2296 4873 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4809 2296 4873 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4809 2210 4873 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4809 2210 4873 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4809 2124 4873 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4809 2124 4873 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4809 2038 4873 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4809 2038 4873 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4809 1952 4873 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4809 1952 4873 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4809 1866 4873 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4809 1866 4873 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4809 1780 4873 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4809 1780 4873 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4728 2640 4792 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4728 2640 4792 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4728 2554 4792 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4728 2554 4792 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4728 2468 4792 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4728 2468 4792 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4728 2382 4792 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4728 2382 4792 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4728 2296 4792 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4728 2296 4792 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4728 2210 4792 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4728 2210 4792 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4728 2124 4792 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4728 2124 4792 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4728 2038 4792 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4728 2038 4792 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4728 1952 4792 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4728 1952 4792 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4728 1866 4792 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4728 1866 4792 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4728 1780 4792 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4728 1780 4792 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4647 2640 4711 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4647 2640 4711 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4647 2554 4711 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4647 2554 4711 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4647 2468 4711 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4647 2468 4711 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4647 2382 4711 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4647 2382 4711 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4647 2296 4711 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4647 2296 4711 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4647 2210 4711 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4647 2210 4711 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4647 2124 4711 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4647 2124 4711 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4647 2038 4711 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4647 2038 4711 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4647 1952 4711 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4647 1952 4711 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4647 1866 4711 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4647 1866 4711 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4647 1780 4711 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4647 1780 4711 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4566 2640 4630 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4566 2640 4630 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4566 2554 4630 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4566 2554 4630 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4566 2468 4630 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4566 2468 4630 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4566 2382 4630 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4566 2382 4630 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4566 2296 4630 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4566 2296 4630 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4566 2210 4630 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4566 2210 4630 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4566 2124 4630 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4566 2124 4630 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4566 2038 4630 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4566 2038 4630 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4566 1952 4630 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4566 1952 4630 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4566 1866 4630 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4566 1866 4630 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4566 1780 4630 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4566 1780 4630 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4485 2640 4549 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4485 2640 4549 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4485 2554 4549 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4485 2554 4549 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4485 2468 4549 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4485 2468 4549 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4485 2382 4549 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4485 2382 4549 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4485 2296 4549 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4485 2296 4549 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4485 2210 4549 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4485 2210 4549 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4485 2124 4549 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4485 2124 4549 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4485 2038 4549 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4485 2038 4549 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4485 1952 4549 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4485 1952 4549 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4485 1866 4549 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4485 1866 4549 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4485 1780 4549 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4485 1780 4549 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4404 2640 4468 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4404 2640 4468 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4404 2554 4468 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4404 2554 4468 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4404 2468 4468 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4404 2468 4468 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4404 2382 4468 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4404 2382 4468 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4404 2296 4468 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4404 2296 4468 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4404 2210 4468 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4404 2210 4468 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4404 2124 4468 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4404 2124 4468 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4404 2038 4468 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4404 2038 4468 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4404 1952 4468 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4404 1952 4468 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4404 1866 4468 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4404 1866 4468 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4404 1780 4468 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4404 1780 4468 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4323 2640 4387 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4323 2640 4387 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4323 2554 4387 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4323 2554 4387 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4323 2468 4387 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4323 2468 4387 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4323 2382 4387 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4323 2382 4387 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4323 2296 4387 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4323 2296 4387 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4323 2210 4387 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4323 2210 4387 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4323 2124 4387 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4323 2124 4387 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4323 2038 4387 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4323 2038 4387 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4323 1952 4387 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4323 1952 4387 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4323 1866 4387 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4323 1866 4387 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4323 1780 4387 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4323 1780 4387 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4242 2640 4306 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4242 2640 4306 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4242 2554 4306 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4242 2554 4306 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4242 2468 4306 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4242 2468 4306 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4242 2382 4306 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4242 2382 4306 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4242 2296 4306 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4242 2296 4306 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4242 2210 4306 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4242 2210 4306 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4242 2124 4306 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4242 2124 4306 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4242 2038 4306 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4242 2038 4306 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4242 1952 4306 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4242 1952 4306 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4242 1866 4306 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4242 1866 4306 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4242 1780 4306 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4242 1780 4306 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4161 2640 4225 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4161 2640 4225 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4161 2554 4225 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4161 2554 4225 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4161 2468 4225 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4161 2468 4225 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4161 2382 4225 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4161 2382 4225 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4161 2296 4225 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4161 2296 4225 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4161 2210 4225 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4161 2210 4225 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4161 2124 4225 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4161 2124 4225 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4161 2038 4225 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4161 2038 4225 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4161 1952 4225 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4161 1952 4225 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4161 1866 4225 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4161 1866 4225 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4161 1780 4225 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4161 1780 4225 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4080 2640 4144 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4080 2640 4144 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4080 2554 4144 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4080 2554 4144 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4080 2468 4144 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4080 2468 4144 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4080 2382 4144 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4080 2382 4144 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4080 2296 4144 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4080 2296 4144 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4080 2210 4144 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4080 2210 4144 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4080 2124 4144 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4080 2124 4144 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4080 2038 4144 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4080 2038 4144 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4080 1952 4144 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4080 1952 4144 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4080 1866 4144 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4080 1866 4144 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 4080 1780 4144 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 4080 1780 4144 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3999 2640 4063 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3999 2640 4063 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3999 2554 4063 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3999 2554 4063 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3999 2468 4063 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3999 2468 4063 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3999 2382 4063 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3999 2382 4063 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3999 2296 4063 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3999 2296 4063 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3999 2210 4063 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3999 2210 4063 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3999 2124 4063 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3999 2124 4063 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3999 2038 4063 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3999 2038 4063 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3999 1952 4063 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3999 1952 4063 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3999 1866 4063 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3999 1866 4063 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3999 1780 4063 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3999 1780 4063 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3918 2640 3982 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3918 2640 3982 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3918 2554 3982 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3918 2554 3982 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3918 2468 3982 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3918 2468 3982 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3918 2382 3982 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3918 2382 3982 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3918 2296 3982 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3918 2296 3982 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3918 2210 3982 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3918 2210 3982 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3918 2124 3982 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3918 2124 3982 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3918 2038 3982 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3918 2038 3982 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3918 1952 3982 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3918 1952 3982 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3918 1866 3982 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3918 1866 3982 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3918 1780 3982 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3918 1780 3982 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3837 2640 3901 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3837 2640 3901 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3837 2554 3901 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3837 2554 3901 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3837 2468 3901 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3837 2468 3901 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3837 2382 3901 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3837 2382 3901 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3837 2296 3901 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3837 2296 3901 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3837 2210 3901 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3837 2210 3901 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3837 2124 3901 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3837 2124 3901 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3837 2038 3901 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3837 2038 3901 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3837 1952 3901 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3837 1952 3901 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3837 1866 3901 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3837 1866 3901 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3837 1780 3901 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3837 1780 3901 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3756 2640 3820 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3756 2640 3820 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3756 2554 3820 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3756 2554 3820 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3756 2468 3820 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3756 2468 3820 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3756 2382 3820 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3756 2382 3820 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3756 2296 3820 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3756 2296 3820 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3756 2210 3820 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3756 2210 3820 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3756 2124 3820 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3756 2124 3820 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3756 2038 3820 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3756 2038 3820 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3756 1952 3820 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3756 1952 3820 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3756 1866 3820 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3756 1866 3820 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3756 1780 3820 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3756 1780 3820 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3675 2640 3739 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3675 2640 3739 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3675 2554 3739 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3675 2554 3739 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3675 2468 3739 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3675 2468 3739 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3675 2382 3739 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3675 2382 3739 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3675 2296 3739 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3675 2296 3739 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3675 2210 3739 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3675 2210 3739 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3675 2124 3739 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3675 2124 3739 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3675 2038 3739 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3675 2038 3739 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3675 1952 3739 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3675 1952 3739 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3675 1866 3739 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3675 1866 3739 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3675 1780 3739 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3675 1780 3739 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3594 2640 3658 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3594 2640 3658 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3594 2554 3658 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3594 2554 3658 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3594 2468 3658 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3594 2468 3658 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3594 2382 3658 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3594 2382 3658 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3594 2296 3658 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3594 2296 3658 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3594 2210 3658 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3594 2210 3658 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3594 2124 3658 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3594 2124 3658 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3594 2038 3658 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3594 2038 3658 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3594 1952 3658 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3594 1952 3658 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3594 1866 3658 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3594 1866 3658 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3594 1780 3658 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3594 1780 3658 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3513 2640 3577 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3513 2640 3577 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3513 2554 3577 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3513 2554 3577 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3513 2468 3577 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3513 2468 3577 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3513 2382 3577 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3513 2382 3577 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3513 2296 3577 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3513 2296 3577 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3513 2210 3577 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3513 2210 3577 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3513 2124 3577 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3513 2124 3577 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3513 2038 3577 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3513 2038 3577 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3513 1952 3577 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3513 1952 3577 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3513 1866 3577 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3513 1866 3577 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3513 1780 3577 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3513 1780 3577 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3432 2640 3496 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3432 2640 3496 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3432 2554 3496 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3432 2554 3496 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3432 2468 3496 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3432 2468 3496 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3432 2382 3496 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3432 2382 3496 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3432 2296 3496 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3432 2296 3496 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3432 2210 3496 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3432 2210 3496 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3432 2124 3496 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3432 2124 3496 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3432 2038 3496 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3432 2038 3496 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3432 1952 3496 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3432 1952 3496 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3432 1866 3496 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3432 1866 3496 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3432 1780 3496 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3432 1780 3496 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3351 2640 3415 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3351 2640 3415 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3351 2554 3415 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3351 2554 3415 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3351 2468 3415 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3351 2468 3415 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3351 2382 3415 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3351 2382 3415 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3351 2296 3415 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3351 2296 3415 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3351 2210 3415 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3351 2210 3415 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3351 2124 3415 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3351 2124 3415 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3351 2038 3415 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3351 2038 3415 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3351 1952 3415 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3351 1952 3415 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3351 1866 3415 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3351 1866 3415 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3351 1780 3415 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3351 1780 3415 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3270 2640 3334 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3270 2640 3334 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3270 2554 3334 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3270 2554 3334 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3270 2468 3334 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3270 2468 3334 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3270 2382 3334 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3270 2382 3334 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3270 2296 3334 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3270 2296 3334 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3270 2210 3334 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3270 2210 3334 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3270 2124 3334 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3270 2124 3334 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3270 2038 3334 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3270 2038 3334 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3270 1952 3334 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3270 1952 3334 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3270 1866 3334 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3270 1866 3334 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3270 1780 3334 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3270 1780 3334 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3189 2640 3253 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3189 2640 3253 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3189 2554 3253 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3189 2554 3253 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3189 2468 3253 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3189 2468 3253 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3189 2382 3253 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3189 2382 3253 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3189 2296 3253 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3189 2296 3253 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3189 2210 3253 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3189 2210 3253 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3189 2124 3253 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3189 2124 3253 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3189 2038 3253 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3189 2038 3253 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3189 1952 3253 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3189 1952 3253 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3189 1866 3253 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3189 1866 3253 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3189 1780 3253 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3189 1780 3253 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3108 2640 3172 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3108 2640 3172 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3108 2554 3172 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3108 2554 3172 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3108 2468 3172 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3108 2468 3172 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3108 2382 3172 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3108 2382 3172 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3108 2296 3172 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3108 2296 3172 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3108 2210 3172 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3108 2210 3172 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3108 2124 3172 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3108 2124 3172 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3108 2038 3172 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3108 2038 3172 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3108 1952 3172 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3108 1952 3172 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3108 1866 3172 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3108 1866 3172 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3108 1780 3172 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3108 1780 3172 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3027 2640 3091 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3027 2640 3091 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3027 2554 3091 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3027 2554 3091 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3027 2468 3091 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3027 2468 3091 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3027 2382 3091 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3027 2382 3091 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3027 2296 3091 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3027 2296 3091 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3027 2210 3091 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3027 2210 3091 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3027 2124 3091 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3027 2124 3091 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3027 2038 3091 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3027 2038 3091 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3027 1952 3091 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3027 1952 3091 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3027 1866 3091 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3027 1866 3091 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 3027 1780 3091 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 3027 1780 3091 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2946 2640 3010 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2946 2640 3010 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2946 2554 3010 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2946 2554 3010 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2946 2468 3010 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2946 2468 3010 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2946 2382 3010 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2946 2382 3010 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2946 2296 3010 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2946 2296 3010 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2946 2210 3010 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2946 2210 3010 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2946 2124 3010 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2946 2124 3010 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2946 2038 3010 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2946 2038 3010 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2946 1952 3010 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2946 1952 3010 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2946 1866 3010 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2946 1866 3010 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2946 1780 3010 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2946 1780 3010 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2865 2640 2929 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2865 2640 2929 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2865 2554 2929 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2865 2554 2929 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2865 2468 2929 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2865 2468 2929 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2865 2382 2929 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2865 2382 2929 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2865 2296 2929 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2865 2296 2929 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2865 2210 2929 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2865 2210 2929 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2865 2124 2929 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2865 2124 2929 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2865 2038 2929 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2865 2038 2929 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2865 1952 2929 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2865 1952 2929 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2865 1866 2929 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2865 1866 2929 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2865 1780 2929 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2865 1780 2929 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2784 2640 2848 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2784 2640 2848 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2784 2554 2848 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2784 2554 2848 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2784 2468 2848 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2784 2468 2848 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2784 2382 2848 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2784 2382 2848 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2784 2296 2848 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2784 2296 2848 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2784 2210 2848 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2784 2210 2848 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2784 2124 2848 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2784 2124 2848 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2784 2038 2848 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2784 2038 2848 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2784 1952 2848 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2784 1952 2848 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2784 1866 2848 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2784 1866 2848 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2784 1780 2848 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2784 1780 2848 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2703 2640 2767 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2703 2640 2767 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2703 2554 2767 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2703 2554 2767 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2703 2468 2767 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2703 2468 2767 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2703 2382 2767 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2703 2382 2767 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2703 2296 2767 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2703 2296 2767 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2703 2210 2767 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2703 2210 2767 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2703 2124 2767 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2703 2124 2767 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2703 2038 2767 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2703 2038 2767 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2703 1952 2767 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2703 1952 2767 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2703 1866 2767 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2703 1866 2767 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2703 1780 2767 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2703 1780 2767 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2622 2640 2686 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2622 2640 2686 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2622 2554 2686 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2622 2554 2686 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2622 2468 2686 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2622 2468 2686 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2622 2382 2686 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2622 2382 2686 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2622 2296 2686 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2622 2296 2686 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2622 2210 2686 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2622 2210 2686 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2622 2124 2686 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2622 2124 2686 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2622 2038 2686 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2622 2038 2686 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2622 1952 2686 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2622 1952 2686 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2622 1866 2686 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2622 1866 2686 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2622 1780 2686 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2622 1780 2686 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2541 2640 2605 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2541 2640 2605 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2541 2554 2605 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2541 2554 2605 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2541 2468 2605 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2541 2468 2605 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2541 2382 2605 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2541 2382 2605 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2541 2296 2605 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2541 2296 2605 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2541 2210 2605 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2541 2210 2605 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2541 2124 2605 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2541 2124 2605 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2541 2038 2605 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2541 2038 2605 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2541 1952 2605 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2541 1952 2605 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2541 1866 2605 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2541 1866 2605 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2541 1780 2605 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2541 1780 2605 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2460 2640 2524 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2460 2640 2524 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2460 2554 2524 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2460 2554 2524 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2460 2468 2524 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2460 2468 2524 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2460 2382 2524 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2460 2382 2524 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2460 2296 2524 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2460 2296 2524 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2460 2210 2524 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2460 2210 2524 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2460 2124 2524 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2460 2124 2524 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2460 2038 2524 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2460 2038 2524 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2460 1952 2524 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2460 1952 2524 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2460 1866 2524 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2460 1866 2524 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2460 1780 2524 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2460 1780 2524 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2379 2640 2443 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2379 2640 2443 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2379 2554 2443 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2379 2554 2443 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2379 2468 2443 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2379 2468 2443 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2379 2382 2443 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2379 2382 2443 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2379 2296 2443 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2379 2296 2443 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2379 2210 2443 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2379 2210 2443 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2379 2124 2443 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2379 2124 2443 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2379 2038 2443 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2379 2038 2443 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2379 1952 2443 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2379 1952 2443 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2379 1866 2443 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2379 1866 2443 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2379 1780 2443 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2379 1780 2443 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2298 2640 2362 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2298 2640 2362 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2298 2554 2362 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2298 2554 2362 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2298 2468 2362 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2298 2468 2362 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2298 2382 2362 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2298 2382 2362 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2298 2296 2362 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2298 2296 2362 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2298 2210 2362 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2298 2210 2362 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2298 2124 2362 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2298 2124 2362 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2298 2038 2362 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2298 2038 2362 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2298 1952 2362 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2298 1952 2362 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2298 1866 2362 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2298 1866 2362 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2298 1780 2362 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2298 1780 2362 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2217 2640 2281 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2217 2640 2281 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2217 2554 2281 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2217 2554 2281 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2217 2468 2281 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2217 2468 2281 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2217 2382 2281 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2217 2382 2281 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2217 2296 2281 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2217 2296 2281 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2217 2210 2281 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2217 2210 2281 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2217 2124 2281 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2217 2124 2281 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2217 2038 2281 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2217 2038 2281 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2217 1952 2281 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2217 1952 2281 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2217 1866 2281 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2217 1866 2281 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2217 1780 2281 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2217 1780 2281 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2136 2640 2200 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2136 2640 2200 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2136 2554 2200 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2136 2554 2200 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2136 2468 2200 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2136 2468 2200 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2136 2382 2200 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2136 2382 2200 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2136 2296 2200 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2136 2296 2200 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2136 2210 2200 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2136 2210 2200 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2136 2124 2200 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2136 2124 2200 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2136 2038 2200 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2136 2038 2200 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2136 1952 2200 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2136 1952 2200 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2136 1866 2200 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2136 1866 2200 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2136 1780 2200 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2136 1780 2200 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2055 2640 2119 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2055 2640 2119 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2055 2554 2119 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2055 2554 2119 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2055 2468 2119 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2055 2468 2119 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2055 2382 2119 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2055 2382 2119 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2055 2296 2119 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2055 2296 2119 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2055 2210 2119 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2055 2210 2119 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2055 2124 2119 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2055 2124 2119 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2055 2038 2119 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2055 2038 2119 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2055 1952 2119 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2055 1952 2119 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2055 1866 2119 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2055 1866 2119 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 2055 1780 2119 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 2055 1780 2119 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1974 2640 2038 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1974 2640 2038 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1974 2554 2038 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1974 2554 2038 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1974 2468 2038 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1974 2468 2038 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1974 2382 2038 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1974 2382 2038 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1974 2296 2038 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1974 2296 2038 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1974 2210 2038 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1974 2210 2038 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1974 2124 2038 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1974 2124 2038 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1974 2038 2038 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1974 2038 2038 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1974 1952 2038 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1974 1952 2038 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1974 1866 2038 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1974 1866 2038 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1974 1780 2038 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1974 1780 2038 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1893 2640 1957 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1893 2640 1957 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1893 2554 1957 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1893 2554 1957 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1893 2468 1957 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1893 2468 1957 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1893 2382 1957 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1893 2382 1957 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1893 2296 1957 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1893 2296 1957 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1893 2210 1957 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1893 2210 1957 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1893 2124 1957 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1893 2124 1957 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1893 2038 1957 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1893 2038 1957 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1893 1952 1957 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1893 1952 1957 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1893 1866 1957 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1893 1866 1957 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1893 1780 1957 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1893 1780 1957 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1812 2640 1876 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1812 2640 1876 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1812 2554 1876 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1812 2554 1876 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1812 2468 1876 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1812 2468 1876 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1812 2382 1876 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1812 2382 1876 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1812 2296 1876 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1812 2296 1876 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1812 2210 1876 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1812 2210 1876 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1812 2124 1876 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1812 2124 1876 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1812 2038 1876 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1812 2038 1876 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1812 1952 1876 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1812 1952 1876 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1812 1866 1876 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1812 1866 1876 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1812 1780 1876 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1812 1780 1876 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1731 2640 1795 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1731 2640 1795 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1731 2554 1795 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1731 2554 1795 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1731 2468 1795 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1731 2468 1795 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1731 2382 1795 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1731 2382 1795 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1731 2296 1795 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1731 2296 1795 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1731 2210 1795 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1731 2210 1795 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1731 2124 1795 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1731 2124 1795 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1731 2038 1795 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1731 2038 1795 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1731 1952 1795 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1731 1952 1795 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1731 1866 1795 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1731 1866 1795 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1731 1780 1795 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1731 1780 1795 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1650 2640 1714 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1650 2640 1714 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1650 2554 1714 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1650 2554 1714 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1650 2468 1714 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1650 2468 1714 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1650 2382 1714 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1650 2382 1714 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1650 2296 1714 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1650 2296 1714 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1650 2210 1714 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1650 2210 1714 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1650 2124 1714 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1650 2124 1714 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1650 2038 1714 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1650 2038 1714 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1650 1952 1714 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1650 1952 1714 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1650 1866 1714 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1650 1866 1714 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1650 1780 1714 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1650 1780 1714 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1569 2640 1633 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1569 2640 1633 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1569 2554 1633 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1569 2554 1633 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1569 2468 1633 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1569 2468 1633 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1569 2382 1633 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1569 2382 1633 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1569 2296 1633 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1569 2296 1633 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1569 2210 1633 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1569 2210 1633 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1569 2124 1633 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1569 2124 1633 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1569 2038 1633 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1569 2038 1633 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1569 1952 1633 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1569 1952 1633 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1569 1866 1633 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1569 1866 1633 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1569 1780 1633 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1569 1780 1633 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1488 2640 1552 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1488 2640 1552 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1488 2554 1552 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1488 2554 1552 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1488 2468 1552 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1488 2468 1552 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1488 2382 1552 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1488 2382 1552 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1488 2296 1552 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1488 2296 1552 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1488 2210 1552 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1488 2210 1552 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1488 2124 1552 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1488 2124 1552 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1488 2038 1552 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1488 2038 1552 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1488 1952 1552 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1488 1952 1552 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1488 1866 1552 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1488 1866 1552 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1488 1780 1552 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1488 1780 1552 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1407 2640 1471 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1407 2640 1471 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1407 2554 1471 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1407 2554 1471 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1407 2468 1471 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1407 2468 1471 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1407 2382 1471 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1407 2382 1471 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1407 2296 1471 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1407 2296 1471 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1407 2210 1471 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1407 2210 1471 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1407 2124 1471 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1407 2124 1471 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1407 2038 1471 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1407 2038 1471 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1407 1952 1471 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1407 1952 1471 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1407 1866 1471 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1407 1866 1471 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1407 1780 1471 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1407 1780 1471 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1326 2640 1390 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1326 2640 1390 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1326 2554 1390 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1326 2554 1390 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1326 2468 1390 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1326 2468 1390 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1326 2382 1390 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1326 2382 1390 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1326 2296 1390 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1326 2296 1390 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1326 2210 1390 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1326 2210 1390 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1326 2124 1390 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1326 2124 1390 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1326 2038 1390 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1326 2038 1390 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1326 1952 1390 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1326 1952 1390 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1326 1866 1390 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1326 1866 1390 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1326 1780 1390 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1326 1780 1390 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1245 2640 1309 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1245 2640 1309 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1245 2554 1309 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1245 2554 1309 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1245 2468 1309 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1245 2468 1309 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1245 2382 1309 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1245 2382 1309 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1245 2296 1309 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1245 2296 1309 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1245 2210 1309 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1245 2210 1309 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1245 2124 1309 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1245 2124 1309 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1245 2038 1309 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1245 2038 1309 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1245 1952 1309 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1245 1952 1309 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1245 1866 1309 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1245 1866 1309 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1245 1780 1309 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1245 1780 1309 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1164 2640 1228 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1164 2640 1228 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1164 2554 1228 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1164 2554 1228 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1164 2468 1228 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1164 2468 1228 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1164 2382 1228 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1164 2382 1228 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1164 2296 1228 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1164 2296 1228 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1164 2210 1228 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1164 2210 1228 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1164 2124 1228 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1164 2124 1228 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1164 2038 1228 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1164 2038 1228 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1164 1952 1228 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1164 1952 1228 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1164 1866 1228 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1164 1866 1228 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1164 1780 1228 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1164 1780 1228 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1083 2640 1147 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1083 2640 1147 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1083 2554 1147 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1083 2554 1147 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1083 2468 1147 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1083 2468 1147 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1083 2382 1147 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1083 2382 1147 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1083 2296 1147 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1083 2296 1147 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1083 2210 1147 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1083 2210 1147 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1083 2124 1147 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1083 2124 1147 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1083 2038 1147 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1083 2038 1147 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1083 1952 1147 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1083 1952 1147 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1083 1866 1147 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1083 1866 1147 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1083 1780 1147 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1083 1780 1147 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1002 2640 1066 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1002 2640 1066 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1002 2554 1066 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1002 2554 1066 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1002 2468 1066 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1002 2468 1066 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1002 2382 1066 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1002 2382 1066 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1002 2296 1066 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1002 2296 1066 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1002 2210 1066 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1002 2210 1066 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1002 2124 1066 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1002 2124 1066 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1002 2038 1066 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1002 2038 1066 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1002 1952 1066 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1002 1952 1066 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1002 1866 1066 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1002 1866 1066 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 1002 1780 1066 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 1002 1780 1066 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 921 2640 985 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 921 2640 985 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 921 2554 985 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 921 2554 985 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 921 2468 985 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 921 2468 985 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 921 2382 985 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 921 2382 985 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 921 2296 985 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 921 2296 985 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 921 2210 985 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 921 2210 985 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 921 2124 985 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 921 2124 985 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 921 2038 985 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 921 2038 985 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 921 1952 985 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 921 1952 985 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 921 1866 985 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 921 1866 985 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 921 1780 985 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 921 1780 985 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 840 2640 904 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 840 2640 904 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 840 2554 904 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 840 2554 904 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 840 2468 904 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 840 2468 904 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 840 2382 904 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 840 2382 904 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 840 2296 904 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 840 2296 904 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 840 2210 904 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 840 2210 904 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 840 2124 904 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 840 2124 904 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 840 2038 904 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 840 2038 904 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 840 1952 904 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 840 1952 904 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 840 1866 904 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 840 1866 904 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 840 1780 904 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 840 1780 904 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 759 2640 823 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 759 2640 823 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 759 2554 823 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 759 2554 823 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 759 2468 823 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 759 2468 823 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 759 2382 823 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 759 2382 823 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 759 2296 823 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 759 2296 823 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 759 2210 823 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 759 2210 823 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 759 2124 823 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 759 2124 823 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 759 2038 823 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 759 2038 823 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 759 1952 823 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 759 1952 823 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 759 1866 823 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 759 1866 823 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 759 1780 823 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 759 1780 823 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 678 2640 742 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 678 2640 742 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 678 2554 742 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 678 2554 742 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 678 2468 742 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 678 2468 742 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 678 2382 742 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 678 2382 742 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 678 2296 742 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 678 2296 742 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 678 2210 742 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 678 2210 742 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 678 2124 742 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 678 2124 742 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 678 2038 742 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 678 2038 742 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 678 1952 742 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 678 1952 742 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 678 1866 742 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 678 1866 742 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 678 1780 742 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 678 1780 742 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 597 2640 661 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 597 2640 661 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 597 2554 661 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 597 2554 661 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 597 2468 661 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 597 2468 661 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 597 2382 661 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 597 2382 661 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 597 2296 661 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 597 2296 661 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 597 2210 661 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 597 2210 661 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 597 2124 661 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 597 2124 661 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 597 2038 661 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 597 2038 661 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 597 1952 661 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 597 1952 661 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 597 1866 661 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 597 1866 661 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 597 1780 661 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 597 1780 661 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 515 2640 579 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 515 2640 579 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 515 2554 579 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 515 2554 579 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 515 2468 579 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 515 2468 579 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 515 2382 579 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 515 2382 579 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 515 2296 579 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 515 2296 579 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 515 2210 579 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 515 2210 579 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 515 2124 579 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 515 2124 579 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 515 2038 579 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 515 2038 579 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 515 1952 579 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 515 1952 579 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 515 1866 579 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 515 1866 579 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 515 1780 579 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 515 1780 579 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 433 2640 497 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 433 2640 497 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 433 2554 497 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 433 2554 497 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 433 2468 497 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 433 2468 497 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 433 2382 497 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 433 2382 497 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 433 2296 497 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 433 2296 497 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 433 2210 497 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 433 2210 497 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 433 2124 497 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 433 2124 497 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 433 2038 497 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 433 2038 497 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 433 1952 497 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 433 1952 497 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 433 1866 497 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 433 1866 497 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 433 1780 497 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 433 1780 497 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 351 2640 415 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 351 2640 415 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 351 2554 415 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 351 2554 415 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 351 2468 415 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 351 2468 415 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 351 2382 415 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 351 2382 415 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 351 2296 415 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 351 2296 415 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 351 2210 415 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 351 2210 415 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 351 2124 415 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 351 2124 415 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 351 2038 415 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 351 2038 415 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 351 1952 415 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 351 1952 415 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 351 1866 415 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 351 1866 415 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 351 1780 415 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 351 1780 415 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 269 2640 333 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 269 2640 333 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 269 2554 333 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 269 2554 333 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 269 2468 333 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 269 2468 333 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 269 2382 333 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 269 2382 333 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 269 2296 333 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 269 2296 333 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 269 2210 333 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 269 2210 333 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 269 2124 333 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 269 2124 333 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 269 2038 333 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 269 2038 333 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 269 1952 333 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 269 1952 333 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 269 1866 333 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 269 1866 333 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal4 s 269 1780 333 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 269 1780 333 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 187 2640 251 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 187 2554 251 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 187 2468 251 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 187 2382 251 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 187 2296 251 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 187 2210 251 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 187 2124 251 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 187 2038 251 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 187 1952 251 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 187 1866 251 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 187 1780 251 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 105 2640 169 2704 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 105 2554 169 2618 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 105 2468 169 2532 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 105 2382 169 2446 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 105 2296 169 2360 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 105 2210 169 2274 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 105 2124 169 2188 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 105 2038 169 2102 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 105 1952 169 2016 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 105 1866 169 1930 6 VCCD
port 8 nsew power bidirectional
rlabel metal3 s 105 1780 169 1844 6 VCCD
port 8 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 9 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 9 nsew power bidirectional
rlabel metal4 s 0 2987 193 3677 6 VDDA
port 9 nsew power bidirectional
rlabel metal4 s 14807 2987 15000 3677 6 VDDA
port 9 nsew power bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 10 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 10 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 10 nsew ground bidirectional
rlabel metal4 s 0 8317 254 9247 6 VSSD
port 10 nsew ground bidirectional
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 12 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 27347506
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 27255970
<< end >>
